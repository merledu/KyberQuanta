`timescale 1ns / 1ps
module tb_encryption;

    // Parameters
    parameter k = 3;
    parameter ELL = 16;
    parameter NUM_COEFFS = 256;
    parameter Q = 3329;

    // Signals for the encryption module
    logic [7:0] pk[1183:0];                 
    logic [ELL-1:0] T_hat_0 [0:NUM_COEFFS-1];
    logic [ELL-1:0] T_hat_1 [0:NUM_COEFFS-1];
    logic [ELL-1:0] T_hat_2 [0:NUM_COEFFS-1];
    logic [255:0] rho_t;
    logic [15:0] A [0:2][0:2][0:255];
    logic [7:0] mess [32-1:0];
    logic clk;
    logic rst;
    logic  done9_mul;
    logic done10_mul;
    logic done11_mul;
                logic [11:0] y [0:2][255:0];
                logic [11:0] e1 [0:2][255:0];
                logic [11:0] e2 [255:0];
                logic [255:0] r;
                logic [15:0] y_ntt [0:2][255:0];
             logic [15:0] mult_out_00 [255:0];
                             logic [15:0] mult_out_01 [255:0];
                             logic [15:0] mult_out_02 [255:0];
                            
                             logic [15:0] mult_out_10 [255:0];
                             logic [15:0] mult_out_11 [255:0];
                             logic [15:0] mult_out_12 [255:0];
                            
                             logic [15:0] mult_out_20 [255:0];
                             logic [15:0] mult_out_21 [255:0];
                             logic [15:0] mult_out_22 [255:0];
                             logic [15:0] mult_out_1 [255:0];
                             logic [15:0] mult_out_2 [255:0];
                             logic [15:0] mult_out_3 [255:0];
                             logic start_mul;           
                             logic  done0_ntt;
                             logic done1_ntt;
                             logic done2_ntt;
                             logic done0_mul;
                               logic  done1_mul;
                                  logic  done2_mul;
                                   logic  done3_mul;
                                   logic  done4_mul;
                                   logic  done5_mul;
                                       logic  done6_mul;
                                     logic done7_mul;
                                     logic  done8_mul;
logic [31:0] in_1 [256-1:0];
logic [31:0] in_2 [256-1:0];
logic [31:0] in_3 [256-1:0];
logic [ 16-1:0] m_dec [0:256-1];
logic start_ntt;
logic start_inverse;
logic done10_ntt;
logic done11_ntt;
logic done12_ntt;
logic [15:0] mul_add [0:2][255:0];
logic [15:0] mul_add_t[0:2][255:0];
logic [31:0] u [0:2][255:0];
logic  [15:0] decom_out [0:256-1];
logic [15:0] result [0:2][255:0];
logic [15:0] com_out [0:2][255:0];
logic [15:0] comp_v [0:2][255:0];
logic [7:0] encode_u [0:2] [320-1:0];
logic [7:0] encode_v [0:2] [320-1:0];

    // Instantiate the encryption module
    encryption #(
        .k(k),
        .ELL(ELL),
        .NUM_COEFFS(NUM_COEFFS),
        .Q(Q)
    ) enc_inst (
    
    .y(y),
    .e1(e1),
    .r(r),
     .e2(e2),
        .pk(pk),
        .T_hat_0(T_hat_0),
        .T_hat_1(T_hat_1),
        .T_hat_2(T_hat_2),
        .rho_t(rho_t),
        .A(A),
        . done9_mul( done9_mul),
        . done10_mul( done10_mul),
        . done11_mul( done11_mul),
                .clk(clk),
                .rst(rst) ,
                 .done0_ntt(done0_ntt),
                 .done1_ntt(done1_ntt),
                .done2_ntt(done2_ntt),
                .mess(mess),
                                                                . mult_out_00( mult_out_00),
                                                                 . mult_out_01( mult_out_01),
                                                                  . mult_out_02( mult_out_02),
                                                                  . mult_out_10( mult_out_10),
                                                                   . mult_out_11( mult_out_11),
                                                                    . mult_out_12( mult_out_12),
                                                                      . mult_out_20( mult_out_20),
                                                                      . mult_out_21( mult_out_21),
                                                                      . mult_out_22( mult_out_22),
                                                                   .y_ntt(y_ntt),
                                                                   .start_ntt(start_ntt),
                                                                   .mult_out_1(mult_out_1),
                                                                   .mult_out_2(mult_out_2),
                                                                   .mult_out_3(mult_out_3),
                                                                     .done0_mul(done0_mul),
                                                                      .done1_mul(done1_mul),
                                                                       .done2_mul(done2_mul),
                                                                        .done3_mul(done3_mul),
                                                                         .done4_mul(done4_mul),
                                                                         .done5_mul(done5_mul),
                                                                         .done6_mul(done6_mul),
                                                                         .done7_mul(done7_mul),
                                                                        .done8_mul(done8_mul),
                                                                        .start_mul(start_mul),  
                                                                        .m_dec(m_dec),    
                                                                   .in_1(in_1),
                                                                   .in_2(in_2),
                                                                   .in_3(in_3),
//                                                                   .u(u),
                                                                   .done10_ntt(done10_ntt),
                                                                   .done11_ntt(done11_ntt),
                                                                   .done12_ntt(done12_ntt),
                                                                   .start_inverse(start_inverse),
                                                                   .mul_add(mul_add),
                                                                   .mul_add_t(mul_add_t),
                                                                   .decom_out(decom_out),
                                                                   .u(u),
                                                                   .result(result),
                                                                   .com_out(com_out),
                                                                   .comp_v(comp_v),
                                                                   .encode_u(encode_u),
                                                                   .encode_v (encode_v )
                                                                   
                                                                   
                                                                  
//                                                                   

//                               .done9_shake(done9_shake)
    );

    // Clock generation
     always begin
           #5 clk = ~clk; // Toggle clock every 5 time units (100 MHz clock)
       end
   
       // Reset and stimulus generation
       initial begin
           // Initialize signals
           clk = 0;
           rst = 0;
       
            pk[0] = 8'ha8;
            pk[1] = 8'he6;
            pk[2] = 8'h51;
            pk[3] = 8'ha1;
            pk[4] = 8'he6;
            pk[5] = 8'h85;
            pk[6] = 8'hf2;
            pk[7] = 8'h24;
            pk[8] = 8'h78;
            pk[9] = 8'ha8;
            pk[10] = 8'h95;
            pk[11] = 8'h4f;
            pk[12] = 8'h00;
            pk[13] = 8'h7b;
            pk[14] = 8'hc7;
            pk[15] = 8'h71;
            pk[16] = 8'h1b;
            pk[17] = 8'h93;
            pk[18] = 8'h07;
            pk[19] = 8'h72;
            pk[20] = 8'hc7;
            pk[21] = 8'h8f;
            pk[22] = 8'h09;
            pk[23] = 8'h2e;
            pk[24] = 8'h82;
            pk[25] = 8'h87;
            pk[26] = 8'h8e;
            pk[27] = 8'h3e;
            pk[28] = 8'h93;
            pk[29] = 8'h7f;
            pk[30] = 8'h36;
            pk[31] = 8'h79;
            pk[32] = 8'h67;
            pk[33] = 8'h53;
            pk[34] = 8'h29;
            pk[35] = 8'h13;
            pk[36] = 8'ha8;
            pk[37] = 8'hd5;
            pk[38] = 8'h3d;
            pk[39] = 8'hfd;
            pk[40] = 8'hf4;
            pk[41] = 8'hbf;
            pk[42] = 8'hb1;
            pk[43] = 8'hf8;
            pk[44] = 8'h84;
            pk[45] = 8'h67;
            pk[46] = 8'h46;
            pk[47] = 8'h59;
            pk[48] = 8'h67;
            pk[49] = 8'h05;
            pk[50] = 8'hcf;
            pk[51] = 8'h34;
            pk[52] = 8'h51;
            pk[53] = 8'h42;
            pk[54] = 8'hb9;
            pk[55] = 8'h72;
            pk[56] = 8'ha3;
            pk[57] = 8'hf1;
            pk[58] = 8'h63;
            pk[59] = 8'h25;
            pk[60] = 8'hc4;
            pk[61] = 8'h0c;
            pk[62] = 8'h29;
            pk[63] = 8'h52;
            pk[64] = 8'ha3;
            pk[65] = 8'h7b;
            pk[66] = 8'h25;
            pk[67] = 8'h89;
            pk[68] = 8'h7e;
            pk[69] = 8'h5e;
            pk[70] = 8'hf3;
            pk[71] = 8'h5f;
            pk[72] = 8'hba;
            pk[73] = 8'heb;
            pk[74] = 8'h73;
            pk[75] = 8'ha4;
            pk[76] = 8'hac;
            pk[77] = 8'hbe;
            pk[78] = 8'hb6;
            pk[79] = 8'ha0;
            pk[80] = 8'hb8;
            pk[81] = 8'h99;
            pk[82] = 8'h42;
            pk[83] = 8'hce;
            pk[84] = 8'hb1;
            pk[85] = 8'h95;
            pk[86] = 8'h53;
            pk[87] = 8'h1c;
            pk[88] = 8'hfc;
            pk[89] = 8'h0a;
            pk[90] = 8'h07;
            pk[91] = 8'h99;
            pk[92] = 8'h39;
            pk[93] = 8'h54;
            pk[94] = 8'h48;
            pk[95] = 8'h3e;
            pk[96] = 8'h6c;
            pk[97] = 8'hbc;
            pk[98] = 8'h87;
            pk[99] = 8'hc0;
            pk[100] = 8'h6a;
            pk[101] = 8'ha7;
            pk[102] = 8'h4f;
            pk[103] = 8'hf0;
            pk[104] = 8'hca;
            pk[105] = 8'hc5;
            pk[106] = 8'h20;
            pk[107] = 8'h7e;
            pk[108] = 8'h53;
            pk[109] = 8'h5b;
            pk[110] = 8'h26;
            pk[111] = 8'h0a;
            pk[112] = 8'ha9;
            pk[113] = 8'h8d;
            pk[114] = 8'h11;
            pk[115] = 8'h98;
            pk[116] = 8'hc0;
            pk[117] = 8'h7d;
            pk[118] = 8'ha6;
            pk[119] = 8'h05;
            pk[120] = 8'hc4;
            pk[121] = 8'hd1;
            pk[122] = 8'h10;
            pk[123] = 8'h20;
            pk[124] = 8'hf6;
            pk[125] = 8'hc9;
            pk[126] = 8'hf7;
            pk[127] = 8'hbb;
            pk[128] = 8'h68;
            pk[129] = 8'hbb;
            pk[130] = 8'h34;
            pk[131] = 8'h56;
            pk[132] = 8'hc7;
            pk[133] = 8'h3a;
            pk[134] = 8'h01;
            pk[135] = 8'hb7;
            pk[136] = 8'h10;
            pk[137] = 8'hbc;
            pk[138] = 8'h99;
            pk[139] = 8'hd1;
            pk[140] = 8'h77;
            pk[141] = 8'h39;
            pk[142] = 8'ha5;
            pk[143] = 8'h17;
            pk[144] = 8'h16;
            pk[145] = 8'haa;
            pk[146] = 8'h01;
            pk[147] = 8'h66;
            pk[148] = 8'h0c;
            pk[149] = 8'h8b;
            pk[150] = 8'h62;
            pk[151] = 8'h8b;
            pk[152] = 8'h2f;
            pk[153] = 8'h56;
            pk[154] = 8'h02;
            pk[155] = 8'hba;
            pk[156] = 8'h65;
            pk[157] = 8'hf0;
            pk[158] = 8'h7e;
            pk[159] = 8'ha9;
            pk[160] = 8'h93;
            pk[161] = 8'h33;
            pk[162] = 8'h6e;
            pk[163] = 8'h89;
            pk[164] = 8'h6e;
            pk[165] = 8'h83;
            pk[166] = 8'hf2;
            pk[167] = 8'hc5;
            pk[168] = 8'h73;
            pk[169] = 8'h1b;
            pk[170] = 8'hbf;
            pk[171] = 8'h03;
            pk[172] = 8'h46;
            pk[173] = 8'h0c;
            pk[174] = 8'h5b;
            pk[175] = 8'h6c;
            pk[176] = 8'h8a;
            pk[177] = 8'hfe;
            pk[178] = 8'hcb;
            pk[179] = 8'h74;
            pk[180] = 8'h8e;
            pk[181] = 8'he3;
            pk[182] = 8'h91;
            pk[183] = 8'he9;
            pk[184] = 8'h89;
            pk[185] = 8'h34;
            pk[186] = 8'ha2;
            pk[187] = 8'hc5;
            pk[188] = 8'h7d;
            pk[189] = 8'h4d;
            pk[190] = 8'h06;
            pk[191] = 8'h9f;
            pk[192] = 8'h50;
            pk[193] = 8'hd8;
            pk[194] = 8'h8b;
            pk[195] = 8'h30;
            pk[196] = 8'hd6;
            pk[197] = 8'h96;
            pk[198] = 8'h6f;
            pk[199] = 8'h38;
            pk[200] = 8'hc3;
            pk[201] = 8'h7b;
            pk[202] = 8'hc6;
            pk[203] = 8'h49;
            pk[204] = 8'hb8;
            pk[205] = 8'h26;
            pk[206] = 8'h34;
            pk[207] = 8'hce;
            pk[208] = 8'h77;
            pk[209] = 8'h22;
            pk[210] = 8'h64;
            pk[211] = 8'h5c;
            pk[212] = 8'hcd;
            pk[213] = 8'h62;
            pk[214] = 8'h50;
            pk[215] = 8'h63;
            pk[216] = 8'h36;
            pk[217] = 8'h46;
            pk[218] = 8'h46;
            pk[219] = 8'hd6;
            pk[220] = 8'hd6;
            pk[221] = 8'h99;
            pk[222] = 8'hdb;
            pk[223] = 8'h57;
            pk[224] = 8'hb4;
            pk[225] = 8'h5e;
            pk[226] = 8'hb6;
            pk[227] = 8'h74;
            pk[228] = 8'h65;
            pk[229] = 8'he1;
            pk[230] = 8'h6d;
            pk[231] = 8'he4;
            pk[232] = 8'hd4;
            pk[233] = 8'h06;
            pk[234] = 8'ha8;
            pk[235] = 8'h18;
            pk[236] = 8'hb9;
            pk[237] = 8'hea;
            pk[238] = 8'he1;
            pk[239] = 8'hca;
            pk[240] = 8'h91;
            pk[241] = 8'h6a;
            pk[242] = 8'h25;
            pk[243] = 8'h94;
            pk[244] = 8'h48;
            pk[245] = 8'h97;
            pk[246] = 8'h08;
            pk[247] = 8'ha4;
            pk[248] = 8'h3c;
            pk[249] = 8'hea;
            pk[250] = 8'h88;
            pk[251] = 8'hb0;
            pk[252] = 8'h2a;
            pk[253] = 8'h4c;
            pk[254] = 8'h03;
            pk[255] = 8'hd0;
            pk[256] = 8'h9b;
            pk[257] = 8'h44;
            pk[258] = 8'h81;
            pk[259] = 8'h5c;
            pk[260] = 8'h97;
            pk[261] = 8'h10;
            pk[262] = 8'h1c;
            pk[263] = 8'haf;
            pk[264] = 8'h50;
            pk[265] = 8'h48;
            pk[266] = 8'hbb;
            pk[267] = 8'hcb;
            pk[268] = 8'h24;
            pk[269] = 8'h7a;
            pk[270] = 8'he2;
            pk[271] = 8'h36;
            pk[272] = 8'h6c;
            pk[273] = 8'hdc;
            pk[274] = 8'h25;
            pk[275] = 8'h4b;
            pk[276] = 8'ha2;
            pk[277] = 8'h21;
            pk[278] = 8'h29;
            pk[279] = 8'hf4;
            pk[280] = 8'h5b;
            pk[281] = 8'h3b;
            pk[282] = 8'h0e;
            pk[283] = 8'hb3;
            pk[284] = 8'h99;
            pk[285] = 8'hca;
            pk[286] = 8'h91;
            pk[287] = 8'ha3;
            pk[288] = 8'h03;
            pk[289] = 8'h40;
            pk[290] = 8'h28;
            pk[291] = 8'h30;
            pk[292] = 8'hec;
            pk[293] = 8'h01;
            pk[294] = 8'hdb;
            pk[295] = 8'h7b;
            pk[296] = 8'h2c;
            pk[297] = 8'ha4;
            pk[298] = 8'h80;
            pk[299] = 8'hcf;
            pk[300] = 8'h35;
            pk[301] = 8'h04;
            pk[302] = 8'h09;
            pk[303] = 8'hb2;
            pk[304] = 8'h16;
            pk[305] = 8'h09;
            pk[306] = 8'h4b;
            pk[307] = 8'h7b;
            pk[308] = 8'h0c;
            pk[309] = 8'h3a;
            pk[310] = 8'he3;
            pk[311] = 8'h3c;
            pk[312] = 8'he1;
            pk[313] = 8'h0a;
            pk[314] = 8'h91;
            pk[315] = 8'h24;
            pk[316] = 8'he8;
            pk[317] = 8'h96;
            pk[318] = 8'h51;
            pk[319] = 8'hab;
            pk[320] = 8'h90;
            pk[321] = 8'h1e;
            pk[322] = 8'ha2;
            pk[323] = 8'h53;
            pk[324] = 8'hc8;
            pk[325] = 8'h41;
            pk[326] = 8'h5b;
            pk[327] = 8'hd7;
            pk[328] = 8'h82;
            pk[329] = 8'h5f;
            pk[330] = 8'h02;
            pk[331] = 8'hbb;
            pk[332] = 8'h22;
            pk[333] = 8'h93;
            pk[334] = 8'h69;
            pk[335] = 8'haf;
            pk[336] = 8'h97;
            pk[337] = 8'h20;
            pk[338] = 8'h28;
            pk[339] = 8'hf2;
            pk[340] = 8'h28;
            pk[341] = 8'h75;
            pk[342] = 8'hea;
            pk[343] = 8'h55;
            pk[344] = 8'haf;
            pk[345] = 8'h16;
            pk[346] = 8'hd3;
            pk[347] = 8'hbc;
            pk[348] = 8'h69;
            pk[349] = 8'hf7;
            pk[350] = 8'h0c;
            pk[351] = 8'h2e;
            pk[352] = 8'he8;
            pk[353] = 8'hb7;
            pk[354] = 8'h5f;
            pk[355] = 8'h28;
            pk[356] = 8'hb4;
            pk[357] = 8'h7d;
            pk[358] = 8'hd3;
            pk[359] = 8'h91;
            pk[360] = 8'hf9;
            pk[361] = 8'h89;
            pk[362] = 8'had;
            pk[363] = 8'he3;
            pk[364] = 8'h14;
            pk[365] = 8'h72;
            pk[366] = 8'h9c;
            pk[367] = 8'h33;
            pk[368] = 8'h1f;
            pk[369] = 8'ha0;
            pk[370] = 8'h4c;
            pk[371] = 8'h19;
            pk[372] = 8'h17;
            pk[373] = 8'hb2;
            pk[374] = 8'h78;
            pk[375] = 8'hc3;
            pk[376] = 8'heb;
            pk[377] = 8'h60;
            pk[378] = 8'h28;
            pk[379] = 8'h68;
            pk[380] = 8'h51;
            pk[381] = 8'h28;
            pk[382] = 8'h21;
            pk[383] = 8'had;
            pk[384] = 8'hc8;
            pk[385] = 8'h25;
            pk[386] = 8'hc6;
            pk[387] = 8'h45;
            pk[388] = 8'h77;
            pk[389] = 8'hce;
            pk[390] = 8'h1e;
            pk[391] = 8'h63;
            pk[392] = 8'hb1;
            pk[393] = 8'hd9;
            pk[394] = 8'h64;
            pk[395] = 8'h4a;
            pk[396] = 8'h61;
            pk[397] = 8'h29;
            pk[398] = 8'h48;
            pk[399] = 8'ha3;
            pk[400] = 8'h48;
            pk[401] = 8'h3c;
            pk[402] = 8'h7f;
            pk[403] = 8'h1b;
            pk[404] = 8'h9a;
            pk[405] = 8'h25;
            pk[406] = 8'h80;
            pk[407] = 8'h00;
            pk[408] = 8'he3;
            pk[409] = 8'h01;
            pk[410] = 8'h96;
            pk[411] = 8'h94;
            pk[412] = 8'h4a;
            pk[413] = 8'h40;
            pk[414] = 8'h36;
            pk[415] = 8'h27;
            pk[416] = 8'h60;
            pk[417] = 8'h9c;
            pk[418] = 8'h76;
            pk[419] = 8'hc7;
            pk[420] = 8'hea;
            pk[421] = 8'h6b;
            pk[422] = 8'h5d;
            pk[423] = 8'he0;
            pk[424] = 8'h17;
            pk[425] = 8'h64;
            pk[426] = 8'hd2;
            pk[427] = 8'h43;
            pk[428] = 8'h79;
            pk[429] = 8'h11;
            pk[430] = 8'h7b;
            pk[431] = 8'h9e;
            pk[432] = 8'ha2;
            pk[433] = 8'h98;
            pk[434] = 8'h48;
            pk[435] = 8'hdc;
            pk[436] = 8'h55;
            pk[437] = 8'h5c;
            pk[438] = 8'h45;
            pk[439] = 8'h4b;
            pk[440] = 8'hce;
            pk[441] = 8'hae;
            pk[442] = 8'h1b;
            pk[443] = 8'ha5;
            pk[444] = 8'hcc;
            pk[445] = 8'h72;
            pk[446] = 8'hc7;
            pk[447] = 8'h4a;
            pk[448] = 8'hb9;
            pk[449] = 8'h6b;
            pk[450] = 8'h9c;
            pk[451] = 8'h91;
            pk[452] = 8'hb9;
            pk[453] = 8'h10;
            pk[454] = 8'hd2;
            pk[455] = 8'h6b;
            pk[456] = 8'h88;
            pk[457] = 8'hb2;
            pk[458] = 8'h56;
            pk[459] = 8'h39;
            pk[460] = 8'hd4;
            pk[461] = 8'h77;
            pk[462] = 8'h8a;
            pk[463] = 8'he2;
            pk[464] = 8'h6c;
            pk[465] = 8'h7c;
            pk[466] = 8'h61;
            pk[467] = 8'h51;
            pk[468] = 8'ha1;
            pk[469] = 8'h9c;
            pk[470] = 8'h6c;
            pk[471] = 8'hd7;
            pk[472] = 8'h93;
            pk[473] = 8'h84;
            pk[474] = 8'h54;
            pk[475] = 8'h37;
            pk[476] = 8'h24;
            pk[477] = 8'h65;
            pk[478] = 8'he4;
            pk[479] = 8'hc5;
            pk[480] = 8'hec;
            pk[481] = 8'h29;
            pk[482] = 8'h24;
            pk[483] = 8'h5a;
            pk[484] = 8'hcb;
            pk[485] = 8'h3d;
            pk[486] = 8'hb5;
            pk[487] = 8'h37;
            pk[488] = 8'h9d;
            pk[489] = 8'he3;
            pk[490] = 8'hda;
            pk[491] = 8'hbf;
            pk[492] = 8'ha6;
            pk[493] = 8'h29;
            pk[494] = 8'ha7;
            pk[495] = 8'hc0;
            pk[496] = 8'h4a;
            pk[497] = 8'h83;
            pk[498] = 8'h53;
            pk[499] = 8'ha8;
            pk[500] = 8'h53;
            pk[501] = 8'h0c;
            pk[502] = 8'h95;
            pk[503] = 8'hac;
            pk[504] = 8'hb7;
            pk[505] = 8'h32;
            pk[506] = 8'hbb;
            pk[507] = 8'h4b;
            pk[508] = 8'hb8;
            pk[509] = 8'h19;
            pk[510] = 8'h32;
            pk[511] = 8'hbb;
            pk[512] = 8'h2c;
            pk[513] = 8'ha7;
            pk[514] = 8'ha8;
            pk[515] = 8'h48;
            pk[516] = 8'hcd;
            pk[517] = 8'h36;
            pk[518] = 8'h68;
            pk[519] = 8'h01;
            pk[520] = 8'h44;
            pk[521] = 8'h4a;
            pk[522] = 8'hbe;
            pk[523] = 8'h23;
            pk[524] = 8'hc8;
            pk[525] = 8'h3b;
            pk[526] = 8'h36;
            pk[527] = 8'h6a;
            pk[528] = 8'h87;
            pk[529] = 8'hd6;
            pk[530] = 8'ha3;
            pk[531] = 8'hcf;
            pk[532] = 8'h36;
            pk[533] = 8'h09;
            pk[534] = 8'h24;
            pk[535] = 8'hc0;
            pk[536] = 8'h02;
            pk[537] = 8'hba;
            pk[538] = 8'he9;
            pk[539] = 8'h0a;
            pk[540] = 8'hf6;
            pk[541] = 8'h5c;
            pk[542] = 8'h48;
            pk[543] = 8'h06;
            pk[544] = 8'h0b;
            pk[545] = 8'h37;
            pk[546] = 8'h52;
            pk[547] = 8'hf2;
            pk[548] = 8'hba;
            pk[549] = 8'hdf;
            pk[550] = 8'h1a;
            pk[551] = 8'hb2;
            pk[552] = 8'h72;
            pk[553] = 8'h20;
            pk[554] = 8'h72;
            pk[555] = 8'h55;
            pk[556] = 8'h4a;
            pk[557] = 8'h50;
            pk[558] = 8'h59;
            pk[559] = 8'h75;
            pk[560] = 8'h35;
            pk[561] = 8'h94;
            pk[562] = 8'he6;
            pk[563] = 8'ha7;
            pk[564] = 8'h02;
            pk[565] = 8'h76;
            pk[566] = 8'h1f;
            pk[567] = 8'hc9;
            pk[568] = 8'h76;
            pk[569] = 8'h84;
            pk[570] = 8'hc8;
            pk[571] = 8'hc4;
            pk[572] = 8'ha7;
            pk[573] = 8'h54;
            pk[574] = 8'h0a;
            pk[575] = 8'h6b;
            pk[576] = 8'h07;
            pk[577] = 8'hfb;
            pk[578] = 8'hc9;
            pk[579] = 8'hde;
            pk[580] = 8'h87;
            pk[581] = 8'hc9;
            pk[582] = 8'h74;
            pk[583] = 8'haa;
            pk[584] = 8'h88;
            pk[585] = 8'h09;
            pk[586] = 8'hd9;
            pk[587] = 8'h28;
            pk[588] = 8'hc7;
            pk[589] = 8'hf4;
            pk[590] = 8'hcb;
            pk[591] = 8'hbf;
            pk[592] = 8'h80;
            pk[593] = 8'h45;
            pk[594] = 8'hae;
            pk[595] = 8'ha5;
            pk[596] = 8'hbc;
            pk[597] = 8'h66;
            pk[598] = 8'h78;
            pk[599] = 8'h25;
            pk[600] = 8'hfd;
            pk[601] = 8'h05;
            pk[602] = 8'ha5;
            pk[603] = 8'h21;
            pk[604] = 8'hf1;
            pk[605] = 8'ha4;
            pk[606] = 8'hbf;
            pk[607] = 8'h53;
            pk[608] = 8'h92;
            pk[609] = 8'h10;
            pk[610] = 8'hc7;
            pk[611] = 8'h11;
            pk[612] = 8'h3b;
            pk[613] = 8'hc3;
            pk[614] = 8'h7b;
            pk[615] = 8'h3e;
            pk[616] = 8'h58;
            pk[617] = 8'hb0;
            pk[618] = 8'hcb;
            pk[619] = 8'hfc;
            pk[620] = 8'h53;
            pk[621] = 8'hc8;
            pk[622] = 8'h41;
            pk[623] = 8'hcb;
            pk[624] = 8'hb0;
            pk[625] = 8'h37;
            pk[626] = 8'h1d;
            pk[627] = 8'he2;
            pk[628] = 8'he5;
            pk[629] = 8'h11;
            pk[630] = 8'hb9;
            pk[631] = 8'h89;
            pk[632] = 8'hcb;
            pk[633] = 8'h7c;
            pk[634] = 8'h70;
            pk[635] = 8'hc0;
            pk[636] = 8'h23;
            pk[637] = 8'h36;
            pk[638] = 8'h6d;
            pk[639] = 8'h78;
            pk[640] = 8'hf9;
            pk[641] = 8'hc3;
            pk[642] = 8'h7e;
            pk[643] = 8'hf0;
            pk[644] = 8'h47;
            pk[645] = 8'hf8;
            pk[646] = 8'h72;
            pk[647] = 8'h0b;
            pk[648] = 8'he1;
            pk[649] = 8'hc7;
            pk[650] = 8'h59;
            pk[651] = 8'ha8;
            pk[652] = 8'hd9;
            pk[653] = 8'h6b;
            pk[654] = 8'h93;
            pk[655] = 8'hf6;
            pk[656] = 8'h5a;
            pk[657] = 8'h94;
            pk[658] = 8'h11;
            pk[659] = 8'h4f;
            pk[660] = 8'hfa;
            pk[661] = 8'hf6;
            pk[662] = 8'h0d;
            pk[663] = 8'h9a;
            pk[664] = 8'h81;
            pk[665] = 8'h79;
            pk[666] = 8'h5e;
            pk[667] = 8'h99;
            pk[668] = 8'h5c;
            pk[669] = 8'h71;
            pk[670] = 8'h15;
            pk[671] = 8'h2a;
            pk[672] = 8'h46;
            pk[673] = 8'h91;
            pk[674] = 8'ha5;
            pk[675] = 8'ha6;
            pk[676] = 8'h02;
            pk[677] = 8'ha9;
            pk[678] = 8'he1;
            pk[679] = 8'hf3;
            pk[680] = 8'h59;
            pk[681] = 8'h9e;
            pk[682] = 8'h37;
            pk[683] = 8'hc7;
            pk[684] = 8'h68;
            pk[685] = 8'hc7;
            pk[686] = 8'hbc;
            pk[687] = 8'h10;
            pk[688] = 8'h89;
            pk[689] = 8'h94;
            pk[690] = 8'hc0;
            pk[691] = 8'h66;
            pk[692] = 8'h9f;
            pk[693] = 8'h3a;
            pk[694] = 8'hdc;
            pk[695] = 8'h95;
            pk[696] = 8'h7d;
            pk[697] = 8'h46;
            pk[698] = 8'hb4;
            pk[699] = 8'hb6;
            pk[700] = 8'h25;
            pk[701] = 8'h69;
            pk[702] = 8'h68;
            pk[703] = 8'he2;
            pk[704] = 8'h90;
            pk[705] = 8'hd7;
            pk[706] = 8'h89;
            pk[707] = 8'h2e;
            pk[708] = 8'ha8;
            pk[709] = 8'h54;
            pk[710] = 8'h64;
            pk[711] = 8'hee;
            pk[712] = 8'h7a;
            pk[713] = 8'h75;
            pk[714] = 8'h0f;
            pk[715] = 8'h39;
            pk[716] = 8'hc5;
            pk[717] = 8'he3;
            pk[718] = 8'h15;
            pk[719] = 8'h2c;
            pk[720] = 8'h2d;
            pk[721] = 8'hfc;
            pk[722] = 8'h56;
            pk[723] = 8'hd8;
            pk[724] = 8'hb0;
            pk[725] = 8'hc9;
            pk[726] = 8'h24;
            pk[727] = 8'hba;
            pk[728] = 8'h8a;
            pk[729] = 8'h95;
            pk[730] = 8'h9a;
            pk[731] = 8'h68;
            pk[732] = 8'h09;
            pk[733] = 8'h65;
            pk[734] = 8'h47;
            pk[735] = 8'hf6;
            pk[736] = 8'h64;
            pk[737] = 8'h23;
            pk[738] = 8'hc8;
            pk[739] = 8'h38;
            pk[740] = 8'h98;
            pk[741] = 8'h2a;
            pk[742] = 8'h57;
            pk[743] = 8'h94;
            pk[744] = 8'hb9;
            pk[745] = 8'he1;
            pk[746] = 8'h53;
            pk[747] = 8'h37;
            pk[748] = 8'h71;
            pk[749] = 8'h33;
            pk[750] = 8'h1a;
            pk[751] = 8'h9a;
            pk[752] = 8'h65;
            pk[753] = 8'h6c;
            pk[754] = 8'h28;
            pk[755] = 8'h82;
            pk[756] = 8'h8b;
            pk[757] = 8'heb;
            pk[758] = 8'h91;
            pk[759] = 8'h26;
            pk[760] = 8'ha6;
            pk[761] = 8'h0e;
            pk[762] = 8'h95;
            pk[763] = 8'he8;
            pk[764] = 8'hc5;
            pk[765] = 8'hd9;
            pk[766] = 8'h06;
            pk[767] = 8'h83;
            pk[768] = 8'h2c;
            pk[769] = 8'h77;
            pk[770] = 8'h10;
            pk[771] = 8'h70;
            pk[772] = 8'h55;
            pk[773] = 8'h76;
            pk[774] = 8'hb1;
            pk[775] = 8'hfb;
            pk[776] = 8'h95;
            pk[777] = 8'h07;
            pk[778] = 8'h26;
            pk[779] = 8'h9d;
            pk[780] = 8'hda;
            pk[781] = 8'hf8;
            pk[782] = 8'hc9;
            pk[783] = 8'h5c;
            pk[784] = 8'he9;
            pk[785] = 8'h71;
            pk[786] = 8'h9b;
            pk[787] = 8'h2c;
            pk[788] = 8'ha8;
            pk[789] = 8'hdd;
            pk[790] = 8'h11;
            pk[791] = 8'h2b;
            pk[792] = 8'he1;
            pk[793] = 8'h0b;
            pk[794] = 8'hcc;
            pk[795] = 8'h9f;
            pk[796] = 8'h4a;
            pk[797] = 8'h37;
            pk[798] = 8'hbd;
            pk[799] = 8'h1b;
            pk[800] = 8'h1e;
            pk[801] = 8'hee;
            pk[802] = 8'hb3;
            pk[803] = 8'h3e;
            pk[804] = 8'hcd;
            pk[805] = 8'ha7;
            pk[806] = 8'h6a;
            pk[807] = 8'he9;
            pk[808] = 8'hf6;
            pk[809] = 8'h9a;
            pk[810] = 8'h5d;
            pk[811] = 8'h4b;
            pk[812] = 8'h29;
            pk[813] = 8'h23;
            pk[814] = 8'ha8;
            pk[815] = 8'h69;
            pk[816] = 8'h57;
            pk[817] = 8'h67;
            pk[818] = 8'h1d;
            pk[819] = 8'h61;
            pk[820] = 8'h93;
            pk[821] = 8'h35;
            pk[822] = 8'hbe;
            pk[823] = 8'h1c;
            pk[824] = 8'h4c;
            pk[825] = 8'h2c;
            pk[826] = 8'h77;
            pk[827] = 8'hce;
            pk[828] = 8'h87;
            pk[829] = 8'hc4;
            pk[830] = 8'h1f;
            pk[831] = 8'h98;
            pk[832] = 8'ha8;
            pk[833] = 8'hcc;
            pk[834] = 8'h46;
            pk[835] = 8'h64;
            pk[836] = 8'h60;
            pk[837] = 8'hfa;
            pk[838] = 8'h30;
            pk[839] = 8'h0a;
            pk[840] = 8'haf;
            pk[841] = 8'h5b;
            pk[842] = 8'h30;
            pk[843] = 8'h1f;
            pk[844] = 8'h0a;
            pk[845] = 8'h1d;
            pk[846] = 8'h09;
            pk[847] = 8'hc8;
            pk[848] = 8'h8e;
            pk[849] = 8'h65;
            pk[850] = 8'hda;
            pk[851] = 8'h4d;
            pk[852] = 8'h8e;
            pk[853] = 8'he6;
            pk[854] = 8'h4f;
            pk[855] = 8'h68;
            pk[856] = 8'hc0;
            pk[857] = 8'h21;
            pk[858] = 8'h89;
            pk[859] = 8'hbb;
            pk[860] = 8'hb3;
            pk[861] = 8'h58;
            pk[862] = 8'h4b;
            pk[863] = 8'haf;
            pk[864] = 8'hf7;
            pk[865] = 8'h16;
            pk[866] = 8'hc8;
            pk[867] = 8'h5d;
            pk[868] = 8'hb6;
            pk[869] = 8'h54;
            pk[870] = 8'h04;
            pk[871] = 8'h8a;
            pk[872] = 8'h00;
            pk[873] = 8'h43;
            pk[874] = 8'h33;
            pk[875] = 8'h48;
            pk[876] = 8'h93;
            pk[877] = 8'h93;
            pk[878] = 8'ha0;
            pk[879] = 8'h74;
            pk[880] = 8'h27;
            pk[881] = 8'hcd;
            pk[882] = 8'h3e;
            pk[883] = 8'h21;
            pk[884] = 8'h7e;
            pk[885] = 8'h6a;
            pk[886] = 8'h34;
            pk[887] = 8'h5f;
            pk[888] = 8'h6c;
            pk[889] = 8'h2c;
            pk[890] = 8'h2b;
            pk[891] = 8'h13;
            pk[892] = 8'hc2;
            pk[893] = 8'h7b;
            pk[894] = 8'h33;
            pk[895] = 8'h72;
            pk[896] = 8'h71;
            pk[897] = 8'hc0;
            pk[898] = 8'hb2;
            pk[899] = 8'h7b;
            pk[900] = 8'h2d;
            pk[901] = 8'hba;
            pk[902] = 8'ha0;
            pk[903] = 8'h0d;
            pk[904] = 8'h23;
            pk[905] = 8'h76;
            pk[906] = 8'h00;
            pk[907] = 8'hb5;
            pk[908] = 8'hb5;
            pk[909] = 8'h94;
            pk[910] = 8'he8;
            pk[911] = 8'hcf;
            pk[912] = 8'h2d;
            pk[913] = 8'hd6;
            pk[914] = 8'h25;
            pk[915] = 8'hea;
            pk[916] = 8'h76;
            pk[917] = 8'hcf;
            pk[918] = 8'h0e;
            pk[919] = 8'hd8;
            pk[920] = 8'h99;
            pk[921] = 8'h12;
            pk[922] = 8'h2c;
            pk[923] = 8'h97;
            pk[924] = 8'h96;
            pk[925] = 8'hb4;
            pk[926] = 8'hb0;
            pk[927] = 8'h18;
            pk[928] = 8'h70;
            pk[929] = 8'h04;
            pk[930] = 8'h25;
            pk[931] = 8'h80;
            pk[932] = 8'h49;
            pk[933] = 8'ha4;
            pk[934] = 8'h77;
            pk[935] = 8'hcd;
            pk[936] = 8'h11;
            pk[937] = 8'hd6;
            pk[938] = 8'h8c;
            pk[939] = 8'h49;
            pk[940] = 8'hb9;
            pk[941] = 8'ha0;
            pk[942] = 8'he7;
            pk[943] = 8'hb0;
            pk[944] = 8'h0b;
            pk[945] = 8'hce;
            pk[946] = 8'h8c;
            pk[947] = 8'hac;
            pk[948] = 8'h78;
            pk[949] = 8'h64;
            pk[950] = 8'hcb;
            pk[951] = 8'hb3;
            pk[952] = 8'h75;
            pk[953] = 8'h14;
            pk[954] = 8'h00;
            pk[955] = 8'h84;
            pk[956] = 8'h74;
            pk[957] = 8'h4c;
            pk[958] = 8'h93;
            pk[959] = 8'h06;
            pk[960] = 8'h26;
            pk[961] = 8'h94;
            pk[962] = 8'hca;
            pk[963] = 8'h79;
            pk[964] = 8'h5c;
            pk[965] = 8'h4f;
            pk[966] = 8'h40;
            pk[967] = 8'he7;
            pk[968] = 8'hac;
            pk[969] = 8'hc9;
            pk[970] = 8'hc5;
            pk[971] = 8'ha1;
            pk[972] = 8'h88;
            pk[973] = 8'h40;
            pk[974] = 8'h72;
            pk[975] = 8'hd8;
            pk[976] = 8'hc3;
            pk[977] = 8'h8d;
            pk[978] = 8'haf;
            pk[979] = 8'hb5;
            pk[980] = 8'h01;
            pk[981] = 8'hee;
            pk[982] = 8'h41;
            pk[983] = 8'h84;
            pk[984] = 8'hdd;
            pk[985] = 8'h5a;
            pk[986] = 8'h81;
            pk[987] = 8'h9e;
            pk[988] = 8'hc2;
            pk[989] = 8'h4e;
            pk[990] = 8'hc1;
            pk[991] = 8'h65;
            pk[992] = 8'h12;
            pk[993] = 8'h61;
            pk[994] = 8'hf9;
            pk[995] = 8'h62;
            pk[996] = 8'hb1;
            pk[997] = 8'h7a;
            pk[998] = 8'h72;
            pk[999] = 8'h15;
            pk[1000] = 8'haa;
            pk[1001] = 8'h4a;
            pk[1002] = 8'h74;
            pk[1003] = 8'h8c;
            pk[1004] = 8'h15;
            pk[1005] = 8'h83;
            pk[1006] = 8'h6c;
            pk[1007] = 8'h38;
            pk[1008] = 8'h91;
            pk[1009] = 8'h37;
            pk[1010] = 8'h67;
            pk[1011] = 8'h82;
            pk[1012] = 8'h04;
            pk[1013] = 8'h83;
            pk[1014] = 8'h8d;
            pk[1015] = 8'h71;
            pk[1016] = 8'h95;
            pk[1017] = 8'ha8;
            pk[1018] = 8'h5b;
            pk[1019] = 8'h4f;
            pk[1020] = 8'h98;
            pk[1021] = 8'ha1;
            pk[1022] = 8'hb5;
            pk[1023] = 8'h74;
            pk[1024] = 8'hc4;
            pk[1025] = 8'hcd;
            pk[1026] = 8'h79;
            pk[1027] = 8'h09;
            pk[1028] = 8'hcd;
            pk[1029] = 8'h1f;
            pk[1030] = 8'h83;
            pk[1031] = 8'h3e;
            pk[1032] = 8'hff;
            pk[1033] = 8'hd1;
            pk[1034] = 8'h48;
            pk[1035] = 8'h55;
            pk[1036] = 8'h43;
            pk[1037] = 8'h22;
            pk[1038] = 8'h9d;
            pk[1039] = 8'h37;
            pk[1040] = 8'h48;
            pk[1041] = 8'hd9;
            pk[1042] = 8'hb5;
            pk[1043] = 8'hcd;
            pk[1044] = 8'h6c;
            pk[1045] = 8'h17;
            pk[1046] = 8'hb9;
            pk[1047] = 8'hb3;
            pk[1048] = 8'hb8;
            pk[1049] = 8'h4a;
            pk[1050] = 8'hef;
            pk[1051] = 8'h8b;
            pk[1052] = 8'hce;
            pk[1053] = 8'h13;
            pk[1054] = 8'he6;
            pk[1055] = 8'h83;
            pk[1056] = 8'h73;
            pk[1057] = 8'h36;
            pk[1058] = 8'h59;
            pk[1059] = 8'hc7;
            pk[1060] = 8'h95;
            pk[1061] = 8'h42;
            pk[1062] = 8'hd6;
            pk[1063] = 8'h15;
            pk[1064] = 8'h78;
            pk[1065] = 8'h2a;
            pk[1066] = 8'h71;
            pk[1067] = 8'hcd;
            pk[1068] = 8'hee;
            pk[1069] = 8'he7;
            pk[1070] = 8'h92;
            pk[1071] = 8'hba;
            pk[1072] = 8'hb5;
            pk[1073] = 8'h1b;
            pk[1074] = 8'hdc;
            pk[1075] = 8'h4b;
            pk[1076] = 8'hbf;
            pk[1077] = 8'he8;
            pk[1078] = 8'h30;
            pk[1079] = 8'h8e;
            pk[1080] = 8'h66;
            pk[1081] = 8'h31;
            pk[1082] = 8'h44;
            pk[1083] = 8'hed;
            pk[1084] = 8'he8;
            pk[1085] = 8'h49;
            pk[1086] = 8'h18;
            pk[1087] = 8'h30;
            pk[1088] = 8'had;
            pk[1089] = 8'h98;
            pk[1090] = 8'hb4;
            pk[1091] = 8'h63;
            pk[1092] = 8'h4f;
            pk[1093] = 8'h64;
            pk[1094] = 8'hab;
            pk[1095] = 8'ha8;
            pk[1096] = 8'hb9;
            pk[1097] = 8'hc0;
            pk[1098] = 8'h42;
            pk[1099] = 8'h27;
            pk[1100] = 8'h26;
            pk[1101] = 8'h53;
            pk[1102] = 8'h92;
            pk[1103] = 8'h0f;
            pk[1104] = 8'h38;
            pk[1105] = 8'h0c;
            pk[1106] = 8'h1a;
            pk[1107] = 8'h17;
            pk[1108] = 8'hca;
            pk[1109] = 8'h87;
            pk[1110] = 8'hce;
            pk[1111] = 8'hd7;
            pk[1112] = 8'haa;
            pk[1113] = 8'hc4;
            pk[1114] = 8'h1c;
            pk[1115] = 8'h82;
            pk[1116] = 8'h88;
            pk[1117] = 8'h87;
            pk[1118] = 8'h93;
            pk[1119] = 8'h18;
            pk[1120] = 8'h1a;
            pk[1121] = 8'h6f;
            pk[1122] = 8'h76;
            pk[1123] = 8'he1;
            pk[1124] = 8'h97;
            pk[1125] = 8'hb7;
            pk[1126] = 8'hb9;
            pk[1127] = 8'h0e;
            pk[1128] = 8'hf9;
            pk[1129] = 8'h09;
            pk[1130] = 8'h43;
            pk[1131] = 8'hbb;
            pk[1132] = 8'h38;
            pk[1133] = 8'h44;
            pk[1134] = 8'h91;
            pk[1135] = 8'h29;
            pk[1136] = 8'h11;
            pk[1137] = 8'hd8;
            pk[1138] = 8'h55;
            pk[1139] = 8'h1e;
            pk[1140] = 8'h54;
            pk[1141] = 8'h66;
            pk[1142] = 8'hc5;
            pk[1143] = 8'h76;
            pk[1144] = 8'h7a;
            pk[1145] = 8'hb0;
            pk[1146] = 8'hbc;
            pk[1147] = 8'h61;
            pk[1148] = 8'ha1;
            pk[1149] = 8'ha3;
            pk[1150] = 8'hf7;
            pk[1151] = 8'h36;
            pk[1152] = 8'h16;
            pk[1153] = 8'h2e;
            pk[1154] = 8'hc0;
            pk[1155] = 8'h98;
            pk[1156] = 8'ha9;
            pk[1157] = 8'h00;
            pk[1158] = 8'hb1;
            pk[1159] = 8'h2d;
            pk[1160] = 8'hd8;
            pk[1161] = 8'hfa;
            pk[1162] = 8'hbb;
            pk[1163] = 8'hfb;
            pk[1164] = 8'h3f;
            pk[1165] = 8'he8;
            pk[1166] = 8'hcb;
            pk[1167] = 8'h1d;
            pk[1168] = 8'hc4;
            pk[1169] = 8'he8;
            pk[1170] = 8'h31;
            pk[1171] = 8'h5f;
            pk[1172] = 8'h2a;
            pk[1173] = 8'hf0;
            pk[1174] = 8'hd3;
            pk[1175] = 8'h2f;
            pk[1176] = 8'h00;
            pk[1177] = 8'h17;
            pk[1178] = 8'hae;
            pk[1179] = 8'h13;
            pk[1180] = 8'h6e;
            pk[1181] = 8'h19;
            pk[1182] = 8'hf0;
            pk[1183] = 8'h28;
            
                mess[0] = 8'hF0;
                mess[1] = 8'h00;
                mess[2] = 8'h0d;
                mess[3] = 8'he5;
                mess[4] = 8'h0f;
                mess[5] = 8'h98;
                mess[6] = 8'h17;
                mess[7] = 8'h23;
                mess[8] = 8'hb8;
                mess[9] = 8'h11;
                mess[10] = 8'h0b;
                mess[11] = 8'h74;
                mess[12] = 8'h4c;
                mess[13] = 8'he4;
                mess[14] = 8'h76;
                mess[15] = 8'h3c;
                mess[16] = 8'hb5;
                mess[17] = 8'hda;
                mess[18] = 8'ha3;
                mess[19] = 8'h22;
                mess[20] = 8'h68;
                mess[21] = 8'hcc;
                mess[22] = 8'hb6;
                mess[23] = 8'h4c;
                mess[24] = 8'hcb;
                mess[25] = 8'h6a;
                mess[26] = 8'h94;
                mess[27] = 8'h5e;
                mess[28] = 8'h9f;
                mess[29] = 8'h98;
                mess[30] = 8'ha2;
                mess[31] = 8'hb5;
         r = 256'hcdf7593486798d29417fecfc7e6fce8dbd073e5f5adb8b2ddaa5667c3f5688f6;
//         message = 276'hF0000de50f981723b8110b744ce4763cb5daa32268ccb64ccb6a945e9f98a2b51e1d7;
        // Continue initializing the rest of the public key...

        // Apply reset signal
        rst = 1;
        #10 rst = 0;  // Reset pulse

        // Wait for the encryption module to complete
        #800000;  // Wait for a while to see the results
//        #1000000;  // Wait for a while to see the results

   // Monitor the results (Display rho_t, A, T_hat_0, T_hat_1, T_hat_2)
       
        
//        for (int i = 0; i < 3; i++) begin
//            for (int j = 0; j < 3; j++) begin
//                for (int k = 0; k < 256; k++) begin
//                    $display("A[%0d][%0d][%0d] = %h", i, j, k, A[i][j][k]);
//                end
//            end
//        end
        
        // Display T_hat values
//        $display("T_hat_0 values:");
//        for (int i = 0; i < NUM_COEFFS; i++) begin
//            $display("T_hat_0[%0d]: %h", i, T_hat_0[i]);
//        end

//        $display("T_hat_1 values:");
//        for (int i = 0; i < NUM_COEFFS; i++) begin
//            $display("T_hat_1[%0d]: %h", i, T_hat_1[i]);
//        end

//        $display("T_hat_2 values:");
//        for (int i = 0; i < NUM_COEFFS; i++) begin
//            $display("T_hat_2[%0d]: %h", i, T_hat_2[i]);
//        end
 // message takes the value of datain (hex value)

    // Debugging message value
//$display("Message (from datain) = %h", message);
// Modify the always_ff block that monitors the changes
     // Debugging datain9 value // Debugging datain value
//              $display("rho_t: %h", rho_t);
// Debugging datain9 value

     
//       $display("Message (datain) = %h", message);
//       $display("Z (xof8) = %h", z);
 // Debugging xof9 value
 
       
//                  $display("done1_shake: %b", done10_shake);
//                  $display("done2_shake: %b", done11_shake);
//                  $display("done3_shake: %b", done12_shake);
//                  $display("done4_shake: %b", done13_shake);
//                  $display("done5_shake: %b", done14_shake);
//   $display("done0_shake: %b", done9_shake); 
//                   $display("done0_cbd: %b", done0_cbd); 
//            $display("done1_cbd: %b", done1_cbd);
//     $display("done2_cbd: %b", done2_cbd);
//                                $display("done3_cbd: %b",done3_cbd);
//                                $display("done4_cbd: %b", done4_cbd);
//                                $display("done5_cbd: %b",done5_cbd);
////         $display("done9_shake: %b", done9_shake);
//$display("r0 = %h", r0);
//$display("r1 = %h", r1);
//$display("r2 = %h", r2);
//$display("r3 = %h", r3);
//$display("r4 = %h", r4);
//$display("r5 = %h", r5);
//        $display("mul_00: f = %h, g = %h, h = %p", A[0][0], y_ntt[0], mult_out_00);
//        $display("mul_01: f = %h, g = %h, h = %p", A[0][1], y_ntt[1], mult_out_01);
//        $display("mul_02: f = %h, g = %h, h = %p", A[0][2], y_ntt[2], mult_out_02);

//        $display("mul_10: f = %h, g = %h, h = %p", A[1][0], y_ntt[0], mult_out_10);
//        $display("mul_11: f = %h, g = %h, h = %p", A[1][1], y_ntt[1], mult_out_11);
//        $display("mul_12: f = %h, g = %h, h = %p", A[1][2], y_ntt[2], mult_out_12);

//        $display("mul_20: f = %h, g = %h, h = %p", A[2][0], y_ntt[0], mult_out_20);
//        $display("mul_21: f = %h, g = %h, h = %p", A[2][1], y_ntt[1], mult_out_21);
//        $display("mul_22: f = %h, g = %h, h = %p", A[2][2], y_ntt[2], mult_out_22);

        $dumpfile("encryption_waveform.vcd");  // Specify the VCD file name
        $dumpvars(0, tb_encryption);  // Dump all variables in the testbench to the VCD file

        // End simulation
        $finish;
    end

endmodule