`timescale 1ns / 1ps

module tb_bytes_to_bits;

    localparam BYTE_COUNT = 384; 
    localparam BIT_COUNT = BYTE_COUNT * 8;

    logic [7:0] B [0:BYTE_COUNT-1]; 
    logic [$clog2(BYTE_COUNT):0] len; 
    logic [BIT_COUNT-1:0] b; 

    bytes_to_bits #(
        .BYTE_COUNT(BYTE_COUNT),
        .BIT_COUNT(BIT_COUNT)
    ) uut (
        .B(B),
        .len(len),
        .b(b)
    );
    logic [7:0] test_data [0:BYTE_COUNT-1]; 
    integer i; 

    initial begin
        $display("Starting Test Case 1...");
        len = 384; 

        for (i = 0; i < BYTE_COUNT; i++) begin
            test_data[i] = (i < 256) ? i : 8'h00; 
        end

//        for (i = 0; i < BYTE_COUNT; i++) begin
//            B[i] = test_data[i];
//        end
B = '{25, 215, 74, 213, 71, 42, 139, 43, 170, 210, 165, 103, 2, 201, 179, 181, 81, 14, 243, 146, 72, 88, 6, 29, 87, 249, 13, 217, 161, 160, 31, 236, 47, 87, 197, 26, 136, 136, 5, 52, 27, 97, 124, 81, 85, 57, 89, 119, 80, 131, 92, 62, 215, 160, 51, 176, 57, 215, 36, 145, 51, 44, 93, 244, 166, 155, 109, 242, 97, 113, 135, 122, 209, 229, 10, 197, 1, 0, 190, 71, 40, 120, 102, 133, 218, 122, 115, 158, 132, 63, 240, 212, 89, 34, 215, 40, 30, 33, 13, 94, 130, 185, 68, 101, 47, 72, 98, 207, 179, 217, 2, 222, 96, 175, 208, 161, 100, 71, 27, 38, 20, 74, 29, 122, 56, 9, 101, 3, 9, 89, 17, 118, 46, 186, 121, 98, 196, 81, 29, 5, 161, 40, 242, 120, 30, 203, 61, 31, 91, 177, 36, 66, 55, 97, 26, 186, 185, 36, 153, 31, 138, 39, 50, 226, 112, 50, 53, 121, 32, 241, 151, 199, 105, 45, 96, 169, 68, 68, 114, 37, 140, 180, 87, 193, 183, 27, 119, 153, 84, 105, 243, 169, 98, 243, 171, 166, 105, 150, 20, 252, 204, 234, 116, 30, 33, 198, 0, 196, 53, 123, 191, 171, 69, 41, 39, 195, 212, 65, 191, 142, 215, 49, 82, 247, 92, 8, 245, 64, 225, 134, 172, 202, 51, 38, 244, 34, 200, 75, 152, 141, 119, 230, 26, 230, 24, 89, 207, 133, 65, 248, 146, 9, 228, 152, 48, 64, 197, 97, 118, 84, 128, 136, 82, 182, 73, 184, 153, 163, 153, 174, 194, 200, 187, 168, 165, 66, 243, 69, 171, 242, 129, 63, 101, 233, 167, 145, 211, 44, 194, 215, 96, 38, 251, 141, 12, 148, 182, 87, 72, 154, 187, 72, 125, 164, 162, 192, 227, 134, 141, 60, 244, 127, 28, 187, 47, 167, 156, 83, 207, 246, 38, 71, 119, 192, 155, 23, 124, 145, 49, 84, 132, 210, 179, 11, 12, 162, 31, 85, 173, 210, 60, 87, 225, 145, 28, 63, 8, 107, 202, 210, 23, 152, 72, 110, 180, 123, 124, 88, 87, 115, 129, 192, 159, 82, 82, 88, 45, 27, 39, 167, 213, 184, 224, 96, 206, 120, 32, 156, 200, 43, 174, 77, 166, 6};
        $display("Input Byte Array:");
        for (i = 0; i < len; i++) begin
            $write("B[%0d] = %h ", i, B[i]);
            if (i % 8 == 7) $display(""); 
        end
        $display("");

        #1; 
        $display("Output Bit Array Length: %0d bits", len * 8);

        $display("Output Bit Array:");
        for (i = 0; i < len * 8; i++) begin
            $write("%b", b[i]);
            if (i % 8 == 7) $write(" "); 
            if (i % 64 == 63) $display(""); 
        end
        $display("");
//        $display("Validating output...");
//        for (i = 0; i < len; i++) begin
//            if (b[i*8 +: 8] !== test_data[i]) begin
//                $fatal("Mismatch at byte %0d: Expected %0h, Got %0h", i, test_data[i], b[i*8 +: 8]);
//            end
//        end
//        $display("Test Case 1 Passed!");

        $finish;
    end

endmodule
