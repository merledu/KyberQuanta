`timescale 1ns / 1ps
module encryption #(
    parameter k = 3,
    parameter ELL = 16,
    parameter NUM_COEFFS = 256,
    parameter Q = 3329
)(
  input logic clk,
  input logic rst,
  input logic [7:0] pk[1183:0],    
//  input [255:0] m,     
  input [255:0] r,     
  output logic [15:0] A [0:2][0:2][0:255],
  output logic [ ELL-1:0] T_hat_0 [0:NUM_COEFFS-1],
  output logic [ ELL-1:0] T_hat_1 [0:NUM_COEFFS-1],
  output logic [ ELL-1:0] T_hat_2 [0:NUM_COEFFS-1],
  output logic [ ELL-1:0] m_dec [0:NUM_COEFFS-1],
  output logic [255:0] rho_t,
  input logic [7:0] m [0:32-1],
  output logic [11:0] y [0:2][255:0],
  output logic [11:0] e1 [0:2][255:0],
  output logic [11:0] e2 [255:0],
  output logic [15:0] y_ntt [0:2][255:0],
  output logic start_ntt,
  output logic [15:0] mult_out_00 [255:0],
  output logic [15:0] mult_out_01 [255:0],
  output logic [15:0] mult_out_02 [255:0],
  output logic [15:0] mult_out_10 [255:0],
  output logic [15:0] mult_out_11 [255:0],
  output logic [15:0] mult_out_12 [255:0],
  output logic [15:0] mult_out_20 [255:0],
  output logic [15:0] mult_out_21 [255:0],
      output logic [15:0] mult_out_22 [255:0],
      output logic  done9_mul,
      output logic  done10_mul,
      output logic  done11_mul,
      output logic [15:0] mult_out_1 [255:0],
      output logic [15:0] mult_out_2 [255:0],
      output logic [15:0] mult_out_3 [255:0],
      output logic [31:0] in_1 [256-1:0],
      output logic [31:0] in_2 [256-1:0],
      output logic [31:0] in_3 [256-1:0],
         output logic [31:0] in_4 [256-1:0],
         output logic [31:0] in_5 [256-1:0],
         output logic [31:0] in_6 [256-1:0],
            output logic [31:0] in_7 [256-1:0],
            output logic [31:0] in_8 [256-1:0],
            output logic [31:0] in_9 [256-1:0],
            output logic [31:0] v_in_1[256-1:0],
             output logic [31:0] v_in_2[256-1:0],
              output logic [31:0] v_in_3 [256-1:0],
            output logic done10_ntt,
               output logic done11_ntt,
               output logic done12_ntt,
               output logic done4_ntt,
               output logic done5_ntt,
               output logic done6_ntt,
               output logic done7_ntt,
               output logic done8_ntt,
               output logic done9_ntt,
               output logic done13_ntt,
               output logic done14_ntt,
               output logic done15_ntt,
               output logic start_inverse,
               output logic [31:0] u_1 [255:0],
               output logic [31:0] u_2 [255:0],
               output logic [31:0] u_3 [255:0],
               output logic [31:0] u_4 [255:0],
               output logic [31:0] u_5 [255:0],
               output logic [31:0] u_6 [255:0],
               output logic [31:0] u_7 [255:0],
               output logic [31:0] u_8 [255:0],
               output logic [31:0] u_9 [255:0],
               output logic [31:0] e2_ext [255:0],
               output logic [31:0] v_1 [255:0],
               output logic [31:0] v_2 [255:0],
               output logic [31:0] v_3 [255:0],
               output logic [15:0] result,
               output logic [15:0] decom_out,
               output logic [15:0] com_out 
      );
    

    logic [7:0] pk_slice0 [0:383];
    logic [7:0] pk_slice1 [0:383];
    logic [7:0] pk_slice2 [0:383];
    logic  done9_shake, done10_shake, done11_shake, done12_shake, done13_shake, done14_shake,done15_shake;
    logic  done0_cbd, done1_cbd, done2_cbd, done3_cbd, done4_cbd, done5_cbd,done6_cbd;
    logic [7:0] parse_array1 [767:0];
    logic [7:0] parse_array2 [767:0];
    logic [7:0] parse_array3 [767:0];
    logic [7:0] parse_array4 [767:0];
    logic [7:0] parse_array5 [767:0];
    logic [7:0] parse_array6 [767:0];
    logic [7:0] parse_array7 [767:0];
    logic [7:0] parse_array8 [767:0];
    logic [7:0] parse_array9 [767:0];
    logic start1;
    logic done0, done1, done2, done3, done4, done5, done6, done7, done8, done9;
    logic done0_shake,done1_shake,done2_shake,done3_shake,done4_shake,done5_shake,done6_shake,done7_shake,done8_shake;
    logic all_shake_done;
    logic [7:0] prf_bytes_0 [127:0];
    logic [7:0] prf_bytes_1 [127:0];
    logic [7:0] prf_bytes_2 [127:0];
    logic [7:0] prf_bytes_3 [127:0];
    logic [7:0] prf_bytes_4 [127:0];
    logic [7:0] prf_bytes_5 [127:0];
    logic [7:0] prf_bytes_6 [127:0];
    logic [1023:0] prf_0, prf_1, prf_2, prf_3, prf_4, prf_5, prf_6;
    logic  start_parse, start_cbd, start_prf;
    logic [15:0] zetas [127:0];
    logic ntt_started;
    logic mul;
    logic [268-1:0] r0;
    logic [268-1:0] r1;
    logic [268-1:0] r2;
    logic [268-1:0] r3;
    logic [268-1:0] r4;
    logic [268-1:0] r5;
    logic done0_mul;
    logic  done1_mul;
    logic  done2_mul;
    logic  done3_mul;
    logic  done4_mul;
    logic  done5_mul;
    logic  done6_mul;
    logic done7_mul;
    logic  done8_mul;

    logic start_mul;
    
    logic  done0_ntt;
    logic done1_ntt;
    logic done2_ntt;
    
    assign pk_slice0 = pk[383:0];
    assign pk_slice1 = pk[767:384];
    assign pk_slice2 = pk[1151:768];
   
assign rho_t = {
           pk[1152], pk[1153], pk[1154], pk[1155],
           pk[1156], pk[1157], pk[1158], pk[1159],
           pk[1160], pk[1161], pk[1162], pk[1163],
           pk[1164], pk[1165], pk[1166], pk[1167],
           pk[1168], pk[1169], pk[1170], pk[1171],
           pk[1172], pk[1173], pk[1174], pk[1175],
           pk[1176], pk[1177], pk[1178], pk[1179],
           pk[1180], pk[1181], pk[1182], pk[1183]
       };


    decode #(.ELL(16), .NUM_COEFFS(256), .BYTE_COUNT(384)) dec0 (
        .byte_array(pk_slice0),
        .len(384),
        .coeffs(T_hat_0)
    );

    decode #(.ELL(16), .NUM_COEFFS(256), .BYTE_COUNT(384)) dec1 (
        .byte_array(pk_slice1),
        .len(384),
        .coeffs(T_hat_1)
    );

    decode #(.ELL(16), .NUM_COEFFS(256), .BYTE_COUNT(384)) dec2 (
        .byte_array(pk_slice2),
        .len(384),
        .coeffs(T_hat_2)
    );
    
     
   
   

        
              //--------------------------XOF 1--------------------------------------
    logic [276-1:0] datain;
    logic [6144-1:0] xof;
    
   assign datain = {4'hF,8'h00, 8'h00,rho_t};
   assign message = datain; 
//   assign done0_shake = 1'b1;
    sponge #(
     .msg_len(276),
     .d_len(6144),
     .capacity(256),
     .r(1600 - 256)
 ) shake1(
        .clk(clk),
        .reset(rst),
        .start(start1),
        .message(datain),
        .z(xof),
        .done(done0_shake)
    );
            
           
           //--------------------------XOF 2--------------------------------------
              logic [276-1:0] datain2;
                   logic [6144-1:0] xof2;
//                  assign message = datain2; 
                   assign datain2 = {4'hF ,8'h00, 8'h02,rho_t};     
                    
                   sponge #(
                    .msg_len(276),
                    .d_len(6144),
                    .capacity(256),
                    .r(1600 - 256)
                ) shake2(
                       .clk(clk),
                       .reset(rst),
                       .start(start1),
                       .message(datain2),
                       .z(xof2),
                       .done(done1_shake)
                   ); 
                    
                 //--------------------------XOF 3--------------------------------------
               logic [276-1:0] datain3;
               logic [6144-1:0] xof3;
//                        assign message = datain3;                           
               assign datain3 = {4'hF , 8'h00, 8'h11,rho_t };      
               sponge #(
                    .msg_len(276),
                     .d_len(6144),
                     .capacity(256),
                     .r(1600 - 256)
                                  ) shake3(
                                        .clk(clk),
                                         .reset(rst),
                                         .start(start1),
                                        .message(datain3),
                                          .z(xof3),
                                           .done(done2_shake)
                                                  );
   
                    // --------------------------XOF 4--------------------------------------
              logic [276-1:0] datain4;
              logic [6144-1:0] xof4;
//                                                            assign message = datain4; 
              assign datain4 = {4'hF ,  8'h01 , 8'h00,rho_t };
              sponge #(
                        .msg_len(276),
                         .d_len(6144),
                         .capacity(256),
                         .r(1600 - 256)
                   ) shake4 (
                              .clk(clk),
                             .reset(rst),
                             .start(start1),
                            .message(datain4),
                             .z(xof4),
                             .done( done3_shake)
                                        );        
                  
                    // --------------------------XOF 5--------------------------------------
                         logic [276-1:0] datain5;
                  logic [6144-1:0] xof5;
//                assign message = datain5; 
            assign datain5 = {4'hF ,  8'h01 , 8'h01,rho_t };
        sponge #(
                      .msg_len(276),
                      .d_len(6144),
                      .capacity(256),
                       .r(1600 - 256)
                                       )
                 shake5 (
                         .clk(clk),
                         .reset(rst),
                         .start(start1),
                         .message(datain5),
                         .z(xof5),
                         .done( done4_shake)
                          );  
                 
                    // --------------------------XOF 6--------------------------------------
                       logic [276-1:0] datain6;
                       logic [6144-1:0] xof6;
//                       assign message = datain6; 
                       assign datain6 = {4'hF ,  8'h1 , 8'h2,rho_t };
                       sponge #(
                       .msg_len(276),
                       .d_len(6144),
                       .capacity(256),
                       .r(1600 - 256)
                       ) shake6 (
                       .clk(clk),
                        .reset(rst),
                        .start(start1),
                        .message(datain6),
                        .z(xof6),
                        .done( done5_shake)
                        );
                  
               // --------------------------XOF 7--------------------------------------
                   logic [276-1:0] datain7;
                   logic [6144-1:0] xof7;
//                    assign message = datain7; 
                   assign datain7 = {4'hF ,  8'h02 , 8'h00,rho_t };
                   sponge #(
                   .msg_len(276),
                   .d_len(6144),
                   .capacity(256),
                   .r(1600 - 256)
                   ) shake7 (
                   .clk(clk),
                   .reset(rst),
                   .start(start1),
                   .message(datain7),
                   .z(xof7),
                   .done( done6_shake)
                    );
   
                    // --------------------------XOF 8--------------------------------------
                     logic [276-1:0] datain8;
                     logic [6144-1:0] xof8;
//                     assign message = datain8; 
                     assign datain8 = {4'hF ,  8'h02 , 8'h01,rho_t };
                      sponge #(
                       .msg_len(276),
                       .d_len(6144),
                       .capacity(256),
                        .r(1600 - 256)
                         ) shake8 (
                          .clk(clk),
                           .reset(rst),
                            .start(start1),
                            .message(datain8),
                            .z(xof8),
                             .done( done7_shake)
                              );
                                                                                                          
                                                                                                          // --------------------------XOF 9--------------------------------------
          logic [276-1:0] datain9;
          logic [6144-1:0] xof9;
//        assign message = datain9; 
          assign datain9 = {4'hF ,  8'h2 , 8'h2,rho_t };
          sponge #(
           .msg_len(276),
           .d_len(6144),
           .capacity(256),
           .r(1600 - 256)
            ) shake9 (
            .clk(clk),
            .reset(rst),
            .start(start1),
            .message(datain9),
            .z(xof9),
            .done( done8_shake)
             );
       parse parse_00 (.clk(clk),.rst(rst),.start(done0_shake),.done(done0), .B(parse_array1), .a(A[0][0]));
       parse parse_01 (.clk(clk),.rst(rst),.start(done1_shake),.done(done1),.B(parse_array2), .a(A[0][1]));
       parse parse_02 (.clk(clk),.rst(rst),.start(done2_shake),.done(done2),.B(parse_array3), .a(A[0][2]));
       
       parse parse_10 (.clk(clk),.rst(rst),.start(done3_shake),.done(done3),.B(parse_array4), .a(A[1][0]));
       parse parse_11 (.clk(clk),.rst(rst),.start(done4_shake),.done(done4),.B(parse_array5), .a(A[1][1]));
       parse parse_12 (.clk(clk),.rst(rst),.start(done4_shake),.done(done5),.B(parse_array6), .a(A[1][2]));
       
       parse parse_20 (.clk(clk),.rst(rst),.start(done4_shake),.done(done6),.B(parse_array7), .a(A[2][0]));
       parse parse_21 (.clk(clk),.rst(rst),.start(done4_shake),.done(done7),.B(parse_array8), .a(A[2][1]));
       parse parse_22 (.clk(clk),.rst(rst),.start(done8_shake),.done(done8),.B(parse_array9), .a(A[2][2]));
       


  always_ff @(posedge clk or posedge rst) begin
           if (rst) begin
           ntt_started <=0;
               all_shake_done <= 0;
               mul <= 0;
//                       start_encode <= 0;
                       start_parse  <= 0;
                       start_cbd    <= 0;
                       start_prf    <= 0;
//                       start_ntt <= 0;
           end else begin
                   start_parse  <= 0;
                   start_cbd    <= 0;
                   start_prf    <= 0;
            start1 <= 1;
           zetas[0] = 17; zetas[1] = 2761; zetas[2] = 583; zetas[3] = 2649; zetas[4] = 1637; zetas[5] = 723; zetas[6] = 2288; zetas[7] = 1100;
                   zetas[8] = 1409; zetas[9] = 2662; zetas[10] = 3281; zetas[11] = 233; zetas[12] = 756; zetas[13] = 2156; zetas[14] = 3015; zetas[15] = 3050;
                   zetas[16] = 1703; zetas[17] = 1651; zetas[18] = 2789; zetas[19] = 1789; zetas[20] = 1847; zetas[21] = 952; zetas[22] = 1461; zetas[23] = 2687;
                   zetas[24] = 939; zetas[25] = 2308; zetas[26] = 2437; zetas[27] = 2388; zetas[28] = 733; zetas[29] = 2337; zetas[30] = 268; zetas[31] = 641;
                   zetas[32] = 1584; zetas[33] = 2298; zetas[34] = 2037; zetas[35] = 3220; zetas[36] = 375; zetas[37] = 2549; zetas[38] = 2090; zetas[39] = 1645;
                   zetas[40] = 1063; zetas[41] = 319; zetas[42] = 2773; zetas[43] = 757; zetas[44] = 2099; zetas[45] = 561; zetas[46] = 2466; zetas[47] = 2594;
                   zetas[48] = 2804; zetas[49] = 1092; zetas[50] = 403; zetas[51] = 1026; zetas[52] = 1143; zetas[53] = 2150; zetas[54] = 2775; zetas[55] = 886;
                   zetas[56] = 1722; zetas[57] = 1212; zetas[58] = 1874; zetas[59] = 1029; zetas[60] = 2110; zetas[61] = 2935; zetas[62] = 885; zetas[63] = 2154;
                   zetas[64] = 289; zetas[65] = 331; zetas[66] = 3253; zetas[67] = 1756; zetas[68] = 1197; zetas[69] = 2304; zetas[70] = 2277; zetas[71] = 2055;
                   zetas[72] = 650; zetas[73] = 1977; zetas[74] = 2513; zetas[75] = 632; zetas[76] = 2865; zetas[77] = 33; zetas[78] = 1320; zetas[79] = 1915;
                   zetas[80] = 2319; zetas[81] = 1435; zetas[82] = 807; zetas[83] = 452; zetas[84] = 1438; zetas[85] = 2868; zetas[86] = 1534; zetas[87] = 2402;
                   zetas[88] = 2647; zetas[89] = 2617; zetas[90] = 1481; zetas[91] = 648; zetas[92] = 2474; zetas[93] = 3110; zetas[94] = 1227; zetas[95] = 910;
                   zetas[96] = 296; zetas[97] = 2447; zetas[98] = 1339; zetas[99] = 1476; zetas[100] = 3046; zetas[101] = 56; zetas[102] = 2240; zetas[103] = 1333;
                   zetas[104] = 1426; zetas[105] = 2094; zetas[106] = 535; zetas[107] = 2882; zetas[108] = 2393; zetas[109] = 2879; zetas[110] = 1974; zetas[111] = 821;
                   zetas[112] = 1062; zetas[113] = 1919; zetas[114] = 193; zetas[115] = 797; zetas[116] = 2786; zetas[117] = 3260; zetas[118] = 569; zetas[119] = 1746;
                   zetas[120] = 2642; zetas[121] = 630; zetas[122] = 1897; zetas[123] = 848; zetas[124] = 2580; zetas[125] = 3289; zetas[126] = 1729; zetas[127] = 3328;
            zetas[17] = 2637;
         
         
          for (int i = 0; i < 768; i = i + 1) begin
                           
                                          parse_array1[i] = xof[(i+1)*8-1 -: 8];
                                           parse_array2[i] = xof2[(i+1)*8-1 -: 8];
                                            parse_array3[i] = xof3[(i+1)*8-1 -: 8];
                                             parse_array4[i] = xof4[(i+1)*8-1 -: 8];
                                              parse_array5[i] = xof5[(i+1)*8-1 -: 8];
                                               parse_array6[i] = xof6[(i+1)*8-1 -: 8];
                                                parse_array7[i] = xof7[(i+1)*8-1 -: 8];
                                                 parse_array8[i] = xof8[(i+1)*8-1 -: 8];
                                                  parse_array9[i] = xof9[(i+1)*8-1 -: 8];
                                             
           end
            if (done0_shake && done1_shake && done2_shake && done3_shake
                             && done6_shake && done7_shake && done8_shake  ) begin
                             start_parse <= 1;
                             start1 <= 0; 
                         end
                         
            if (done0 && done1 && done2 && done3 && done4 && done5 && done6 && done7 && done8 && !done9_shake && !done10_shake && !done11_shake && !done12_shake && !done13_shake && !done14_shake) begin
                                                      start_parse <= 0;
                                                      start_prf <= 1;
                                                       
                                                  end
  for (int i = 0; i < 128; i++) begin
                             prf_bytes_0[i] = prf_0[8*i +: 8];
                             prf_bytes_1[i] = prf_1[8*i +: 8];
                             prf_bytes_2[i] = prf_2[8*i +: 8];
                             prf_bytes_3[i] = prf_3[8*i +: 8];
                             prf_bytes_4[i] = prf_4[8*i +: 8];
                             prf_bytes_5[i] = prf_5[8*i +: 8];
                             prf_bytes_6[i] = prf_6[8*i +: 8];
                         end
//            
                  if (done0_shake && done1_shake && done2_shake && done3_shake &&
                      done4_shake && done5_shake && done6_shake && done7_shake && done8_shake) begin
                      all_shake_done <= 1;
                      start1 <= 0; 
                  end else begin
                      all_shake_done <= 0; 
                  end
             
                         
              end
          end
         
     
//     //-----------------prf0-------------------------
    
     
     assign r0 = {4'h1111, 8'h00,r}; 
     assign r1 = {4'h1111, 8'h01,r};
      assign r2 = {4'h1111, 8'h02,r};
         assign r3 = {4'h1111, 8'h03,r};  
            assign r4 = {4'h1111, 8'h04,r}; 
             assign r5 = {4'h1111, 8'h05,r};
             
     sponge #(.msg_len(268),
      .d_len(1024), 
      .capacity(512),
       .r(1600 - 512))
        prf0 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r0),
         .z(prf_0),
         .done(done9_shake)
     );
     
  
     sponge #(.msg_len(268), 
     .d_len(1024), 
     .capacity(512), 
     .r(1600 - 512)) 
     prf1 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r1),
         .z(prf_1),
         .done(done10_shake)
     );
     
    
     sponge #(.msg_len(268), 
     .d_len(1024), 
     .capacity(512),
      .r(1600 - 512)) 
      prf2 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r2),
         .z(prf_2),
         .done(done11_shake)
     );
   
  
     sponge #(.msg_len(268),
      .d_len(1024), 
      .capacity(512),
       .r(1600 - 512))
        prf3 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r3),
         .z(prf_3),
         .done(done12_shake)
     );
     
   
     sponge #(.msg_len(268),
      .d_len(1024),
       .capacity(512),
        .r(1600 - 512)) 
        prf4 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r4),
         .z(prf_4),
         .done(done13_shake)
     );
     
     
    
     sponge #(.msg_len(268),
      .d_len(1024),
       .capacity(512),
        .r(1600 - 512))
      prf5 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r5),
         .z(prf_5),
         .done(done14_shake)
     );
                  
        CBD cbd0 (.clk(clk), .reset(rst), .start(done14_shake), .done(done0_cbd), .byte_array(prf_bytes_0), .len(128), .f(y[0]));
        CBD cbd1 (.clk(clk), .reset(rst), .start(done14_shake), .done(done1_cbd), .byte_array(prf_bytes_1), .len(128), .f(y[1]));
        CBD cbd2 (.clk(clk), .reset(rst), .start(done14_shake), .done(done2_cbd), .byte_array(prf_bytes_2), .len(128), .f(y[2]));
        
        CBD cbd3 (.clk(clk), .reset(rst), .start(done14_shake), .done(done3_cbd), .byte_array(prf_bytes_3), .len(128), .f(e1[0]));
        CBD cbd4 (.clk(clk), .reset(rst), .start(done14_shake), .done(done4_cbd), .byte_array(prf_bytes_4), .len(128), .f(e1[1]));
        CBD cbd5 (.clk(clk), .reset(rst), .start(done14_shake), .done(done5_cbd), .byte_array(prf_bytes_5), .len(128), .f(e1[2]));
        

        logic [268-1:0] r6;
        assign r6 = {4'h1111, 8'h06,r}; 
        sponge #(.msg_len(268),
             .d_len(1024), 
             .capacity(512),
              .r(1600 - 512))
               prf6 (
                .clk(clk),
                .reset(rst),
                .start(done8),
                .message(r6),
                .z(prf_6),
                .done(done15_shake)
            );
               CBD cbd6  (
                  .clk(clk), 
                           .reset(rst), 
                           .start(done14_shake), 
                           .done(done6_cbd), 
                           .byte_array(prf_bytes_6), 
                           .len(128), 
                           .f(e2)
              );
              
               assign start_ntt = (done5_cbd && !done0_ntt && !done1_ntt && !done2_ntt);
               
                   ntt ntt_y0 (.clk(clk), .reset(rst), .f(y[0]), .start(start_ntt), .done(done0_ntt), .f_hat(y_ntt[0]));
                   ntt ntt_y1 (.clk(clk), .reset(rst), .f(y[1]), .start(start_ntt), .done(done1_ntt),.f_hat(y_ntt[1]));
                   ntt ntt_y2 (.clk(clk), .reset(rst), .f(y[2]), .start(start_ntt), .done(done2_ntt),.f_hat(y_ntt[2]));
      
                      multiply_ntts mul_20 (.clk(clk), .reset(rst),.f(A[2][0]), .g(y_ntt[0]),.zetas(zetas), .h(mult_out_20), .start(start_mul),.done(done6_mul));
                      multiply_ntts mul_21 (.clk(clk), .reset(rst),.f(A[2][1]), .g(y_ntt[1]), .zetas(zetas),.h(mult_out_21), .start(start_mul), .done(done7_mul));
                      multiply_ntts mul_22 (.clk(clk), .reset(rst),.f(A[2][2]), .g(y_ntt[2]), .zetas(zetas),.h(mult_out_22), .start(start_mul), .done(done8_mul));
                                           mul_add[0][0] <= ((mult_out_00[0] + mult_out_01[0] + mult_out_02[0])%3329);
                      mul_add[0][1] <= ((mult_out_00[1] + mult_out_01[1] + mult_out_02[1])%3329) ;
                                                                              mul_add[0][2] <= ((mult_out_00[2] + mult_out_01[2] + mult_out_02[2])%3329) ;
                                                                              mul_add[0][3] <= ((mult_out_00[3] + mult_out_01[3] + mult_out_02[3])%3329) ;
                                                                              mul_add[0][4] <= ((mult_out_00[4] + mult_out_01[4] + mult_out_02[4])%3329) ;
                                                                              mul_add[0][5]<=((mult_out_00[5] + mult_out_01[5] + mult_out_02[5])%3329) ;
                                                                              mul_add[0][6]<=((mult_out_00[6] + mult_out_01[6] + mult_out_02[6])%3329);
                                                                              mul_add[0][7]<=((mult_out_00[7] + mult_out_01[7] + mult_out_02[7])%3329) ;
                                                                              mul_add[0][8]<=((mult_out_00[8] + mult_out_01[8] + mult_out_02[8])%3329);
                                                                              mul_add[0][9]<=((mult_out_00[9] + mult_out_01[9] + mult_out_02[9])%3329) ;
                                                                              mul_add[0][10]<=((mult_out_00[10] + mult_out_01[10] + mult_out_02[10])%3329) ;
                                                                              mul_add[0][11]<=((mult_out_00[11] + mult_out_01[11] + mult_out_02[11])%3329) ;
                                                                              mul_add[0][12]<=((mult_out_00[12] + mult_out_01[12] + mult_out_02[12])%3329) ;
                                                                              mul_add[0][13]<=((mult_out_00[13] + mult_out_01[13] + mult_out_02[13])%3329) ;
                                                                              mul_add[0][14]<=((mult_out_00[14] + mult_out_01[14] + mult_out_02[14])%3329) ;
                                                                              mul_add[0][15]<=((mult_out_00[15] + mult_out_01[15] + mult_out_02[15])%3329) ;
                                                                              mul_add[0][16]<=((mult_out_00[16] + mult_out_01[16] + mult_out_02[16])%3329) ;
                                                                              mul_add[0][17]<=((mult_out_00[17] + mult_out_01[17] + mult_out_02[17])%3329) ;
                                                                              mul_add[0][18]<=((mult_out_00[18] + mult_out_01[18] + mult_out_02[18])%3329) ;
                                                                              mul_add[0][19]<=((mult_out_00[19] + mult_out_01[19] + mult_out_02[19])%3329) ;
                                                                              mul_add[0][20]<=((mult_out_00[20] + mult_out_01[20] + mult_out_02[20])%3329) ;
                                                                              mul_add[0][21]<=((mult_out_00[21] + mult_out_01[21] + mult_out_02[21])%3329) ;
                                                                              mul_add[0][22]<=((mult_out_00[22] + mult_out_01[22] + mult_out_02[22])%3329) ;
                                                                              mul_add[0][23]<=((mult_out_00[23] + mult_out_01[23] + mult_out_02[23])%3329) ;
                                                                              mul_add[0][24]<=((mult_out_00[24] + mult_out_01[24] + mult_out_02[24])%3329) ;
                                                                              mul_add[0][25]<=((mult_out_00[25] + mult_out_01[25] + mult_out_02[25])%3329) ;
                                                                              mul_add[0][26]<=((mult_out_00[26] + mult_out_01[26] + mult_out_02[26])%3329) ;
                                                                              mul_add[0][27]<=((mult_out_00[27] + mult_out_01[27] + mult_out_02[27])%3329) ;
                                                                              mul_add[0][28]<=((mult_out_00[28] + mult_out_01[28] + mult_out_02[28])%3329) ;
                                                                              mul_add[0][29]<=((mult_out_00[29] + mult_out_01[29] + mult_out_02[29])%3329) ;
                                                                              mul_add[0][30]<=((mult_out_00[30] + mult_out_01[30] + mult_out_02[30])%3329) ;
                                                                              mul_add[0][31]<=((mult_out_00[31] + mult_out_01[31] + mult_out_02[31])%3329) ;
                                                                              mul_add[0][32]<=((mult_out_00[32] + mult_out_01[32] + mult_out_02[32])%3329) ;
                                                                              mul_add[0][33]<=((mult_out_00[33] + mult_out_01[33] + mult_out_02[33])%3329) ;
                                                                              mul_add[0][34]<=((mult_out_00[34] + mult_out_01[34] + mult_out_02[34])%3329) ;
                                                                              mul_add[0][35]<=((mult_out_00[35] + mult_out_01[35] + mult_out_02[35])%3329) ;
                                                                              mul_add[0][36]<=((mult_out_00[36] + mult_out_01[36] + mult_out_02[36])%3329) ;
                                                                              mul_add[0][37]<=((mult_out_00[37] + mult_out_01[37] + mult_out_02[37])%3329) ;
                                                                              mul_add[0][38]<=((mult_out_00[38] + mult_out_01[38] + mult_out_02[38])%3329) ;
                                                                              mul_add[0][39]<=((mult_out_00[39] + mult_out_01[39] + mult_out_02[39])%3329) ;
                                                                              mul_add[0][40]<=((mult_out_00[40] + mult_out_01[40] + mult_out_02[40])%3329) ;
                                                                              mul_add[0][41]<=((mult_out_00[41] + mult_out_01[41] + mult_out_02[41])%3329) ;
                                                                              mul_add[0][42]<=((mult_out_00[42] + mult_out_01[42] + mult_out_02[42])%3329) ;
                                                                              mul_add[0][43]<=((mult_out_00[43] + mult_out_01[43] + mult_out_02[43])%3329) ;
                                                                              mul_add[0][44]<=((mult_out_00[44] + mult_out_01[44] + mult_out_02[44])%3329) ;
                                                                              mul_add[0][45]<=((mult_out_00[45] + mult_out_01[45] + mult_out_02[45])%3329) ;
                                                                              mul_add[0][46]<=((mult_out_00[46] + mult_out_01[46] + mult_out_02[46])%3329) ;
                                                                              mul_add[0][47]<=((mult_out_00[47] + mult_out_01[47] + mult_out_02[47])%3329) ;
                                                                              mul_add[0][48]<=((mult_out_00[48] + mult_out_01[48] + mult_out_02[48])%3329) ;
                                                                              mul_add[0][49]<=((mult_out_00[49] + mult_out_01[49] + mult_out_02[49])%3329) ;
                                                                              mul_add[0][50]<=((mult_out_00[50] + mult_out_01[50] + mult_out_02[50])%3329) ;
                                                                              mul_add[0][51]<=((mult_out_00[51] + mult_out_01[51] + mult_out_02[51])%3329) ;
                                                                              mul_add[0][52]<=((mult_out_00[52] + mult_out_01[52] + mult_out_02[52])%3329) ;
                                                                              mul_add[0][53]<=((mult_out_00[53] + mult_out_01[53] + mult_out_02[53])%3329) ;
                                                                              mul_add[0][54]<=((mult_out_00[54] + mult_out_01[54] + mult_out_02[54])%3329) ;
                                                                              mul_add[0][55]<=((mult_out_00[55] + mult_out_01[55] + mult_out_02[55])%3329) ;
                                                                              mul_add[0][56]<=((mult_out_00[56] + mult_out_01[56] + mult_out_02[56])%3329) ;
                                                                              mul_add[0][57]<=((mult_out_00[57] + mult_out_01[57] + mult_out_02[57])%3329) ;
                                                                              mul_add[0][58]<=((mult_out_00[58] + mult_out_01[58] + mult_out_02[58])%3329) ;
                                                                              mul_add[0][59]<=((mult_out_00[59] + mult_out_01[59] + mult_out_02[59])%3329) ;
                                                                              mul_add[0][60]<=((mult_out_00[60] + mult_out_01[60] + mult_out_02[60])%3329) ;
                                                                              mul_add[0][61]<=((mult_out_00[61] + mult_out_01[61] + mult_out_02[61])%3329) ;
                                                                              mul_add[0][62]<=((mult_out_00[62] + mult_out_01[62] + mult_out_02[62])%3329) ;
                                                                              mul_add[0][63]<=((mult_out_00[63] + mult_out_01[63] + mult_out_02[63])%3329) ;
                                                                              mul_add[0][64]<=((mult_out_00[64] + mult_out_01[64] + mult_out_02[64])%3329) ;
                                                                              mul_add[0][65]<=((mult_out_00[65] + mult_out_01[65] + mult_out_02[65])%3329) ;
                                                                              mul_add[0][66]<=((mult_out_00[66] + mult_out_01[66] + mult_out_02[66])%3329) ;
                                                                              mul_add[0][67]<=((mult_out_00[67] + mult_out_01[67] + mult_out_02[67])%3329) ;
                                                                              mul_add[0][68]<=((mult_out_00[68] + mult_out_01[68] + mult_out_02[68])%3329) ;
                                                                              mul_add[0][69]<=((mult_out_00[69] + mult_out_01[69] + mult_out_02[69])%3329) ;
                                                                              mul_add[0][70]<=((mult_out_00[70] + mult_out_01[70] + mult_out_02[70])%3329) ;
                                                                              mul_add[0][71]<=((mult_out_00[71] + mult_out_01[71] + mult_out_02[71])%3329) ;
                                                                              mul_add[0][72]<=((mult_out_00[72] + mult_out_01[72] + mult_out_02[72])%3329) ;
                                                                              mul_add[0][73]<=((mult_out_00[73] + mult_out_01[73] + mult_out_02[73])%3329) ;
                                                                              mul_add[0][74]<=((mult_out_00[74] + mult_out_01[74] + mult_out_02[74])%3329) ;
                                                                              mul_add[0][75]<=((mult_out_00[75] + mult_out_01[75] + mult_out_02[75])%3329) ;
                                                                              mul_add[0][76]<=((mult_out_00[76] + mult_out_01[76] + mult_out_02[76])%3329) ;
                                                                              mul_add[0][77]<=((mult_out_00[77] + mult_out_01[77] + mult_out_02[77])%3329) ;
                                                                              mul_add[0][78]<=((mult_out_00[78] + mult_out_01[78] + mult_out_02[78])%3329) ;
                                                                              mul_add[0][79]<=((mult_out_00[79] + mult_out_01[79] + mult_out_02[79])%3329) ;
                                                                              mul_add[0][80]<=((mult_out_00[80] + mult_out_01[80] + mult_out_02[80])%3329) ;
                                                                              mul_add[0][81]<=((mult_out_00[81] + mult_out_01[81] + mult_out_02[81])%3329) ;
                                                                              mul_add[0][82]<=((mult_out_00[82] + mult_out_01[82] + mult_out_02[82])%3329) ;
                                                                              mul_add[0][83]<=((mult_out_00[83] + mult_out_01[83] + mult_out_02[83])%3329) ;
                                                                              mul_add[0][84]<=((mult_out_00[84] + mult_out_01[84] + mult_out_02[84])%3329) ;
                                                                              mul_add[0][85]<=((mult_out_00[85] + mult_out_01[85] + mult_out_02[85])%3329) ;
                                                                              mul_add[0][86]<=((mult_out_00[86] + mult_out_01[86] + mult_out_02[86])%3329) ;
                                                                              mul_add[0][87]<=((mult_out_00[87] + mult_out_01[87] + mult_out_02[87])%3329) ;
                                                                              mul_add[0][88]<=((mult_out_00[88] + mult_out_01[88] + mult_out_02[88])%3329) ;
                                                                              mul_add[0][89]<=((mult_out_00[89] + mult_out_01[89] + mult_out_02[89])%3329) ;
                                                                              mul_add[0][90]<=((mult_out_00[90] + mult_out_01[90] + mult_out_02[90])%3329) ;
                                                                              mul_add[0][91]<=((mult_out_00[91] + mult_out_01[91] + mult_out_02[91])%3329) ;
                                                                              mul_add[0][92]<=((mult_out_00[92] + mult_out_01[92] + mult_out_02[92])%3329) ;
                                                                              mul_add[0][93]<=((mult_out_00[93] + mult_out_01[93] + mult_out_02[93])%3329) ;
                                                                              mul_add[0][94]<=((mult_out_00[94] + mult_out_01[94] + mult_out_02[94])%3329) ;
                                                                              mul_add[0][95]<=((mult_out_00[95] + mult_out_01[95] + mult_out_02[95])%3329) ;
                                                                              mul_add[0][96]<=((mult_out_00[96] + mult_out_01[96] + mult_out_02[96])%3329) ;
                                                                              mul_add[0][97]<=((mult_out_00[97] + mult_out_01[97] + mult_out_02[97])%3329) ;
                                                                              mul_add[0][98]<=((mult_out_00[98] + mult_out_01[98] + mult_out_02[98])%3329) ;
                                                                              mul_add[0][99]<=((mult_out_00[99] + mult_out_01[99] + mult_out_02[99])%3329) ;
                                                                              mul_add[0][100]<=((mult_out_00[100] + mult_out_01[100] + mult_out_02[100])%3329) ;
                                                                              mul_add[0][101]<=((mult_out_00[101] + mult_out_01[101] + mult_out_02[101])%3329) ;
                                                                              mul_add[0][102]<=((mult_out_00[102] + mult_out_01[102] + mult_out_02[102])%3329) ;
                                                                              mul_add[0][103]<=((mult_out_00[103] + mult_out_01[103] + mult_out_02[103])%3329) ;
                                                                              mul_add[0][104]<=((mult_out_00[104] + mult_out_01[104] + mult_out_02[104])%3329) ;
                                                                              mul_add[0][105]<=((mult_out_00[105] + mult_out_01[105] + mult_out_02[105])%3329) ;
                                                                              mul_add[0][106]<=((mult_out_00[106] + mult_out_01[106] + mult_out_02[106])%3329) ;
                                                                              mul_add[0][107]<=((mult_out_00[107] + mult_out_01[107] + mult_out_02[107])%3329) ;
                                                                              mul_add[0][108]<=((mult_out_00[108] + mult_out_01[108] + mult_out_02[108])%3329) ;
                                                                              mul_add[0][109]<=((mult_out_00[109] + mult_out_01[109] + mult_out_02[109])%3329) ;
                                                                              mul_add[0][110]<=((mult_out_00[110] + mult_out_01[110] + mult_out_02[110])%3329) ;
                                                                              mul_add[0][111]<=((mult_out_00[111] + mult_out_01[111] + mult_out_02[111])%3329) ;
                                                                              mul_add[0][112]<=((mult_out_00[112] + mult_out_01[112] + mult_out_02[112])%3329) ;
                                                                              mul_add[0][113]<=((mult_out_00[113] + mult_out_01[113] + mult_out_02[113])%3329) ;
                                                                              mul_add[0][114]<=((mult_out_00[114] + mult_out_01[114] + mult_out_02[114])%3329) ;
                                                                              mul_add[0][115]<=((mult_out_00[115] + mult_out_01[115] + mult_out_02[115])%3329) ;
                                                                              mul_add[0][116]<=((mult_out_00[116] + mult_out_01[116] + mult_out_02[116])%3329) ;
                                                                              mul_add[0][117]<=((mult_out_00[117] + mult_out_01[117] + mult_out_02[117])%3329) ;
                                                                              mul_add[0][118]<=((mult_out_00[118] + mult_out_01[118] + mult_out_02[118])%3329) ;
                                                                              mul_add[0][119]<=((mult_out_00[119] + mult_out_01[119] + mult_out_02[119])%3329) ;
                                                                              mul_add[0][120]<=((mult_out_00[120] + mult_out_01[120] + mult_out_02[120])%3329) ;
                                                                              mul_add[0][121]<=((mult_out_00[121] + mult_out_01[121] + mult_out_02[121])%3329) ;
                                                                              mul_add[0][122]<=((mult_out_00[122] + mult_out_01[122] + mult_out_02[122])%3329) ;
                                                                              mul_add[0][123]<=((mult_out_00[123] + mult_out_01[123] + mult_out_02[123])%3329) ;
                                                                              mul_add[0][124]<=((mult_out_00[124] + mult_out_01[124] + mult_out_02[124])%3329) ;
                                                                              mul_add[0][125]<=((mult_out_00[125] + mult_out_01[125] + mult_out_02[125])%3329) ;
                                                                              mul_add[0][126]<=((mult_out_00[126] + mult_out_01[126] + mult_out_02[126])%3329) ;
                                                                              mul_add[0][127]<=((mult_out_00[127] + mult_out_01[127] + mult_out_02[127])%3329) ;
                                                                              mul_add[0][128]<=((mult_out_00[128] + mult_out_01[128] + mult_out_02[128])%3329) ;
                                                                              mul_add[0][129]<=((mult_out_00[129] + mult_out_01[129] + mult_out_02[129])%3329) ;
                                                                              mul_add[0][130]<=((mult_out_00[130] + mult_out_01[130] + mult_out_02[130])%3329) ;
                                                                              mul_add[0][131]<=((mult_out_00[131] + mult_out_01[131] + mult_out_02[131])%3329) ;
                                                                              mul_add[0][132]<=((mult_out_00[132] + mult_out_01[132] + mult_out_02[132])%3329) ;
                                                                              mul_add[0][133]<=((mult_out_00[133] + mult_out_01[133] + mult_out_02[133])%3329) ;
                                                                              mul_add[0][134]<=((mult_out_00[134] + mult_out_01[134] + mult_out_02[134])%3329) ;
                                                                              mul_add[0][135]<=((mult_out_00[135] + mult_out_01[135] + mult_out_02[135])%3329) ;
                                                                              mul_add[0][136]<=((mult_out_00[136] + mult_out_01[136] + mult_out_02[136])%3329) ;
                                                                              mul_add[0][137]<=((mult_out_00[137] + mult_out_01[137] + mult_out_02[137])%3329) ;
                                                                              mul_add[0][138]<=((mult_out_00[138] + mult_out_01[138] + mult_out_02[138])%3329) ;
                                                                              mul_add[0][139]<=((mult_out_00[139] + mult_out_01[139] + mult_out_02[139])%3329) ;
                                                                              mul_add[0][140]<=((mult_out_00[140] + mult_out_01[140] + mult_out_02[140])%3329) ;
                                                                              mul_add[0][141]<=((mult_out_00[141] + mult_out_01[141] + mult_out_02[141])%3329) ;
                                                                              mul_add[0][142]<=((mult_out_00[142] + mult_out_01[142] + mult_out_02[142])%3329) ;
                                                                              mul_add[0][143]<=((mult_out_00[143] + mult_out_01[143] + mult_out_02[143])%3329) ;
                                                                              mul_add[0][144]<=((mult_out_00[144] + mult_out_01[144] + mult_out_02[144])%3329) ;
                                                                              mul_add[0][145]<=((mult_out_00[145] + mult_out_01[145] + mult_out_02[145])%3329) ;
                                                                              mul_add[0][146]<=((mult_out_00[146] + mult_out_01[146] + mult_out_02[146])%3329) ;
                                                                              mul_add[0][147]<=((mult_out_00[147] + mult_out_01[147] + mult_out_02[147])%3329) ;
                                                                              mul_add[0][148]<=((mult_out_00[148] + mult_out_01[148] + mult_out_02[148])%3329) ;
                                                                              mul_add[0][149]<=((mult_out_00[149] + mult_out_01[149] + mult_out_02[149])%3329) ;
                                                                              mul_add[0][150]<=((mult_out_00[150] + mult_out_01[150] + mult_out_02[150])%3329) ;
                                                                              mul_add[0][151]<=((mult_out_00[151] + mult_out_01[151] + mult_out_02[151])%3329) ;
                                                                              mul_add[0][152]<=((mult_out_00[152] + mult_out_01[152] + mult_out_02[152])%3329) ;
                                                                              mul_add[0][153]<=((mult_out_00[153] + mult_out_01[153] + mult_out_02[153])%3329) ;
                                                                              mul_add[0][154]<=((mult_out_00[154] + mult_out_01[154] + mult_out_02[154])%3329) ;
                                                                              mul_add[0][155]<=((mult_out_00[155] + mult_out_01[155] + mult_out_02[155])%3329) ;
                                                                              mul_add[0][156]<=((mult_out_00[156] + mult_out_01[156] + mult_out_02[156])%3329) ;
                                                                              mul_add[0][157]<=((mult_out_00[157] + mult_out_01[157] + mult_out_02[157])%3329) ;
                                                                              mul_add[0][158]<=((mult_out_00[158] + mult_out_01[158] + mult_out_02[158])%3329) ;
                                                                              mul_add[0][159]<=((mult_out_00[159] + mult_out_01[159] + mult_out_02[159])%3329) ;
                                                                              mul_add[0][160]<=((mult_out_00[160] + mult_out_01[160] + mult_out_02[160])%3329) ;
                                                                              mul_add[0][161]<=((mult_out_00[161] + mult_out_01[161] + mult_out_02[161])%3329) ;
                                                                              mul_add[0][162]<=((mult_out_00[162] + mult_out_01[162] + mult_out_02[162])%3329) ;
                                                                              mul_add[0][163]<=((mult_out_00[163] + mult_out_01[163] + mult_out_02[163])%3329) ;
                                                                              mul_add[0][164]<=((mult_out_00[164] + mult_out_01[164] + mult_out_02[164])%3329) ;
                                                                              mul_add[0][165]<=((mult_out_00[165] + mult_out_01[165] + mult_out_02[165])%3329) ;
                                                                              mul_add[0][166]<=((mult_out_00[166] + mult_out_01[166] + mult_out_02[166])%3329) ;
                                                                              mul_add[0][167]<=((mult_out_00[167] + mult_out_01[167] + mult_out_02[167])%3329) ;
                                                                              mul_add[0][168]<=((mult_out_00[168] + mult_out_01[168] + mult_out_02[168])%3329) ;
                                                                              mul_add[0][169]<=((mult_out_00[169] + mult_out_01[169] + mult_out_02[169])%3329) ;
                                                                              mul_add[0][170]<=((mult_out_00[170] + mult_out_01[170] + mult_out_02[170])%3329) ;
                                                                              mul_add[0][171]<=((mult_out_00[171] + mult_out_01[171] + mult_out_02[171])%3329) ;
                                                                              mul_add[0][172]<=((mult_out_00[172] + mult_out_01[172] + mult_out_02[172])%3329) ;
                                                                              mul_add[0][173]<=((mult_out_00[173] + mult_out_01[173] + mult_out_02[173])%3329) ;
                                                                              mul_add[0][174]<=((mult_out_00[174] + mult_out_01[174] + mult_out_02[174])%3329) ;
                                                                              mul_add[0][175]<=((mult_out_00[175] + mult_out_01[175] + mult_out_02[175])%3329) ;
                                                                              mul_add[0][176]<=((mult_out_00[176] + mult_out_01[176] + mult_out_02[176])%3329) ;
                                                                              mul_add[0][177]<=((mult_out_00[177] + mult_out_01[177] + mult_out_02[177])%3329) ;
                                                                              mul_add[0][178]<=((mult_out_00[178] + mult_out_01[178] + mult_out_02[178])%3329) ;
                                                                              mul_add[0][179]<=((mult_out_00[179] + mult_out_01[179] + mult_out_02[179])%3329) ;
                                                                              mul_add[0][180]<=((mult_out_00[180] + mult_out_01[180] + mult_out_02[180])%3329) ;
                                                                              mul_add[0][181]<=((mult_out_00[181] + mult_out_01[181] + mult_out_02[181])%3329) ;
                                                                              mul_add[0][182]<=((mult_out_00[182] + mult_out_01[182] + mult_out_02[182])%3329) ;
                                                                              mul_add[0][183]<=((mult_out_00[183] + mult_out_01[183] + mult_out_02[183])%3329) ;
                                                                              mul_add[0][184]<=((mult_out_00[184] + mult_out_01[184] + mult_out_02[184])%3329) ;
                                                                              mul_add[0][185]<=((mult_out_00[185] + mult_out_01[185] + mult_out_02[185])%3329) ;
                                                                              mul_add[0][186]<=((mult_out_00[186] + mult_out_01[186] + mult_out_02[186])%3329) ;
                                                                              mul_add[0][187]<=((mult_out_00[187] + mult_out_01[187] + mult_out_02[187])%3329) ;
                                                                              mul_add[0][188]<=((mult_out_00[188] + mult_out_01[188] + mult_out_02[188])%3329) ;
                                                                              mul_add[0][189]<=((mult_out_00[189] + mult_out_01[189] + mult_out_02[189])%3329) ;
                                                                              mul_add[0][190]<=((mult_out_00[190] + mult_out_01[190] + mult_out_02[190])%3329) ;
                                                                              mul_add[0][191]<=((mult_out_00[191] + mult_out_01[191] + mult_out_02[191])%3329) ;
                                                                              mul_add[0][192]<=((mult_out_00[192] + mult_out_01[192] + mult_out_02[192])%3329) ;
                                                                              mul_add[0][193]<=((mult_out_00[193] + mult_out_01[193] + mult_out_02[193])%3329) ;
                                                                              mul_add[0][194]<=((mult_out_00[194] + mult_out_01[194] + mult_out_02[194])%3329) ;
                                                                              mul_add[0][195]<=((mult_out_00[195] + mult_out_01[195] + mult_out_02[195])%3329) ;
                                                                              mul_add[0][196]<=((mult_out_00[196] + mult_out_01[196] + mult_out_02[196])%3329) ;
                                                                              mul_add[0][197]<=((mult_out_00[197] + mult_out_01[197] + mult_out_02[197])%3329) ;
                                                                              mul_add[0][198]<=((mult_out_00[198] + mult_out_01[198] + mult_out_02[198])%3329) ;
                                                                              mul_add[0][199]<=((mult_out_00[199] + mult_out_01[199] + mult_out_02[199])%3329) ;
                                                                              mul_add[0][200]<=((mult_out_00[200] + mult_out_01[200] + mult_out_02[200])%3329) ;
                                                                              mul_add[0][201]<=((mult_out_00[201] + mult_out_01[201] + mult_out_02[201])%3329) ;
                                                                              mul_add[0][202]<=((mult_out_00[202] + mult_out_01[202] + mult_out_02[202])%3329) ;
                                                                              mul_add[0][203]<=((mult_out_00[203] + mult_out_01[203] + mult_out_02[203])%3329) ;
                                                                              mul_add[0][204]<=((mult_out_00[204] + mult_out_01[204] + mult_out_02[204])%3329) ;
                                                                              mul_add[0][205]<=((mult_out_00[205] + mult_out_01[205] + mult_out_02[205])%3329) ;
                                                                              mul_add[0][206]<=((mult_out_00[206] + mult_out_01[206] + mult_out_02[206])%3329) ;
                                                                              mul_add[0][207]<=((mult_out_00[207] + mult_out_01[207] + mult_out_02[207])%3329) ;
                                                                              mul_add[0][208]<=((mult_out_00[208] + mult_out_01[208] + mult_out_02[208])%3329) ;
                                                                              mul_add[0][209]<=((mult_out_00[209] + mult_out_01[209] + mult_out_02[209])%3329) ;
                                                                              mul_add[0][210]<=((mult_out_00[210] + mult_out_01[210] + mult_out_02[210])%3329) ;
                                                                              mul_add[0][211]<=((mult_out_00[211] + mult_out_01[211] + mult_out_02[211])%3329) ;
                                                                              mul_add[0][212]<=((mult_out_00[212] + mult_out_01[212] + mult_out_02[212])%3329) ;
                                                                              mul_add[0][213]<=((mult_out_00[213] + mult_out_01[213] + mult_out_02[213])%3329) ;
                                                                              mul_add[0][214]<=((mult_out_00[214] + mult_out_01[214] + mult_out_02[214])%3329) ;
                                                                              mul_add[0][215]<=((mult_out_00[215] + mult_out_01[215] + mult_out_02[215])%3329) ;
                                                                              mul_add[0][216]<=((mult_out_00[216] + mult_out_01[216] + mult_out_02[216])%3329) ;
                                                                              mul_add[0][217]<=((mult_out_00[217] + mult_out_01[217] + mult_out_02[217])%3329) ;
                                                                              mul_add[0][218]<=((mult_out_00[218] + mult_out_01[218] + mult_out_02[218])%3329) ;
                                                                              mul_add[0][219]<=((mult_out_00[219] + mult_out_01[219] + mult_out_02[219])%3329) ;
                                                                              mul_add[0][220]<=((mult_out_00[220] + mult_out_01[220] + mult_out_02[220])%3329) ;
                                                                              mul_add[0][221]<=((mult_out_00[221] + mult_out_01[221] + mult_out_02[221])%3329) ;
                                                                              mul_add[0][222]<=((mult_out_00[222] + mult_out_01[222] + mult_out_02[222])%3329) ;
                                                                              mul_add[0][223]<=((mult_out_00[223] + mult_out_01[223] + mult_out_02[223])%3329) ;
                                                                              mul_add[0][224]<=((mult_out_00[224] + mult_out_01[224] + mult_out_02[224])%3329) ;
                                                                              mul_add[0][225]<=((mult_out_00[225] + mult_out_01[225] + mult_out_02[225])%3329) ;
                                                                              mul_add[0][226]<=((mult_out_00[226] + mult_out_01[226] + mult_out_02[226])%3329) ;
                                                                              mul_add[0][227]<=((mult_out_00[227] + mult_out_01[227] + mult_out_02[227])%3329) ;
                                                                              mul_add[0][228]<=((mult_out_00[228] + mult_out_01[228] + mult_out_02[228])%3329) ;
                                                                              mul_add[0][229]<=((mult_out_00[229] + mult_out_01[229] + mult_out_02[229])%3329) ;
                                                                              mul_add[0][230]<=((mult_out_00[230] + mult_out_01[230] + mult_out_02[230])%3329) ;
                                                                              mul_add[0][231]<=((mult_out_00[231] + mult_out_01[231] + mult_out_02[231])%3329) ;
                                                                              mul_add[0][232]<=((mult_out_00[232] + mult_out_01[232] + mult_out_02[232])%3329) ;
                                                                              mul_add[0][233]<=((mult_out_00[233] + mult_out_01[233] + mult_out_02[233])%3329) ;
                                                                              mul_add[0][234]<=((mult_out_00[234] + mult_out_01[234] + mult_out_02[234])%3329) ;
                                                                              mul_add[0][235]<=((mult_out_00[235] + mult_out_01[235] + mult_out_02[235])%3329) ;
                                                                              mul_add[0][236]<=((mult_out_00[236] + mult_out_01[236] + mult_out_02[236])%3329) ;
                                                                              mul_add[0][237]<=((mult_out_00[237] + mult_out_01[237] + mult_out_02[237])%3329) ;
                                                                              mul_add[0][238]<=((mult_out_00[238] + mult_out_01[238] + mult_out_02[238])%3329) ;
                                                                              mul_add[0][239]<=((mult_out_00[239] + mult_out_01[239] + mult_out_02[239])%3329) ;
                                                                              mul_add[0][240]<=((mult_out_00[240] + mult_out_01[240] + mult_out_02[240])%3329) ;
                                                                              mul_add[0][241]<=((mult_out_00[241] + mult_out_01[241] + mult_out_02[241])%3329) ;
                                                                              mul_add[0][242]<=((mult_out_00[242] + mult_out_01[242] + mult_out_02[242])%3329) ;
                                                                              mul_add[0][243]<=((mult_out_00[243] + mult_out_01[243] + mult_out_02[243])%3329) ;
                                                                              mul_add[0][244]<=((mult_out_00[244] + mult_out_01[244] + mult_out_02[244])%3329) ;
                                                                              mul_add[0][245]<=((mult_out_00[245] + mult_out_01[245] + mult_out_02[245])%3329) ;
                                                                              mul_add[0][246]<=((mult_out_00[246] + mult_out_01[246] + mult_out_02[246])%3329) ;
                                                                              mul_add[0][247]<=((mult_out_00[247] + mult_out_01[247] + mult_out_02[247])%3329) ;
                                                                              mul_add[0][248]<=((mult_out_00[248] + mult_out_01[248] + mult_out_02[248])%3329) ;
                                                                              mul_add[0][249]<=((mult_out_00[249] + mult_out_01[249] + mult_out_02[249])%3329) ;
                                                                              mul_add[0][250]<=((mult_out_00[250] + mult_out_01[250] + mult_out_02[250])%3329) ;
                                                                              mul_add[0][251]<=((mult_out_00[251] + mult_out_01[251] + mult_out_02[251])%3329) ;
                                                                              mul_add[0][252]<=((mult_out_00[252] + mult_out_01[252] + mult_out_02[252])%3329) ;
                                                                              mul_add[0][253]<=((mult_out_00[253] + mult_out_01[253] + mult_out_02[253])%3329) ;
                                                                              mul_add[0][254]<=((mult_out_00[254] + mult_out_01[254] + mult_out_02[254])%3329) ;
                                                                              mul_add[0][255]<=((mult_out_00[255] + mult_out_01[255] + mult_out_02[255])%3329) ;
                                                                             
                                                                              mul_add[1][0]<=((mult_out_10[0] + mult_out_11[0] + mult_out_12[0])%3329) ;
                                                                              mul_add[1][1]<=((mult_out_10[1] + mult_out_11[1] + mult_out_12[1])%3329) ;
                                                                              mul_add[1][2]<=((mult_out_10[2] + mult_out_11[2] + mult_out_12[2])%3329) ;
                                                                              mul_add[1][3]<=((mult_out_10[3] + mult_out_11[3] + mult_out_12[3])%3329) ;
                                                                              mul_add[1][4]<=((mult_out_10[4] + mult_out_11[4] + mult_out_12[4])%3329) ;
                                                                              mul_add[1][5]<=((mult_out_10[5] + mult_out_11[5] + mult_out_12[5])%3329) ;
                                                                              mul_add[1][6]<=((mult_out_10[6] + mult_out_11[6] + mult_out_12[6])%3329) ;
                                                                              mul_add[1][7]<=((mult_out_10[7] + mult_out_11[7] + mult_out_12[7])%3329) ;
                                                                              mul_add[1][8]<=((mult_out_10[8] + mult_out_11[8] + mult_out_12[8])%3329) ;
                                                                              mul_add[1][9]<=((mult_out_10[9] + mult_out_11[9] + mult_out_12[9])%3329) ;
                                                                              mul_add[1][10]<=((mult_out_10[10] + mult_out_11[10] + mult_out_12[10])%3329) ;
                                                                              mul_add[1][11]<=((mult_out_10[11] + mult_out_11[11] + mult_out_12[11])%3329) ;
                                                                              mul_add[1][12]<=((mult_out_10[12] + mult_out_11[12] + mult_out_12[12])%3329) ;
                                                                              mul_add[1][13]<=((mult_out_10[13] + mult_out_11[13] + mult_out_12[13])%3329) ;
                                                                              mul_add[1][14]<=((mult_out_10[14] + mult_out_11[14] + mult_out_12[14])%3329) ;
                                                                              mul_add[1][15]<=((mult_out_10[15] + mult_out_11[15] + mult_out_12[15])%3329) ;
                                                                              mul_add[1][16]<=((mult_out_10[16] + mult_out_11[16] + mult_out_12[16])%3329) ;
                                                                              mul_add[1][17]<=((mult_out_10[17] + mult_out_11[17] + mult_out_12[17])%3329) ;
                                                                              mul_add[1][18]<=((mult_out_10[18] + mult_out_11[18] + mult_out_12[18])%3329) ;
                                                                              mul_add[1][19]<=((mult_out_10[19] + mult_out_11[19] + mult_out_12[19])%3329) ;
                                                                              mul_add[1][20]<=((mult_out_10[20] + mult_out_11[20] + mult_out_12[20])%3329) ;
                                                                              mul_add[1][21]<=((mult_out_10[21] + mult_out_11[21] + mult_out_12[21])%3329) ;
                                                                              mul_add[1][22]<=((mult_out_10[22] + mult_out_11[22] + mult_out_12[22])%3329) ;
                                                                              mul_add[1][23]<=((mult_out_10[23] + mult_out_11[23] + mult_out_12[23])%3329) ;
                                                                              mul_add[1][24]<=((mult_out_10[24] + mult_out_11[24] + mult_out_12[24])%3329) ;
                                                                              mul_add[1][25]<=((mult_out_10[25] + mult_out_11[25] + mult_out_12[25])%3329) ;
                                                                              mul_add[1][26]<=((mult_out_10[26] + mult_out_11[26] + mult_out_12[26])%3329) ;
                                                                              mul_add[1][27]<=((mult_out_10[27] + mult_out_11[27] + mult_out_12[27])%3329) ;
                                                                              mul_add[1][28]<=((mult_out_10[28] + mult_out_11[28] + mult_out_12[28])%3329) ;
                                                                              mul_add[1][29]<=((mult_out_10[29] + mult_out_11[29] + mult_out_12[29])%3329) ;
                                                                              mul_add[1][30]<=((mult_out_10[30] + mult_out_11[30] + mult_out_12[30])%3329) ;
                                                                              mul_add[1][31]<=((mult_out_10[31] + mult_out_11[31] + mult_out_12[31])%3329) ;
                                                                              mul_add[1][32]<=((mult_out_10[32] + mult_out_11[32] + mult_out_12[32])%3329) ;
                                                                              mul_add[1][33]<=((mult_out_10[33] + mult_out_11[33] + mult_out_12[33])%3329) ;
                                                                              mul_add[1][34]<=((mult_out_10[34] + mult_out_11[34] + mult_out_12[34])%3329) ;
                                                                              mul_add[1][35]<=((mult_out_10[35] + mult_out_11[35] + mult_out_12[35])%3329) ;
                                                                              mul_add[1][36]<=((mult_out_10[36] + mult_out_11[36] + mult_out_12[36])%3329) ;
                                                                              mul_add[1][37]<=((mult_out_10[37] + mult_out_11[37] + mult_out_12[37])%3329) ;
                                                                              mul_add[1][38]<=((mult_out_10[38] + mult_out_11[38] + mult_out_12[38])%3329) ;
                                                                              mul_add[1][39]<=((mult_out_10[39] + mult_out_11[39] + mult_out_12[39])%3329) ;
                                                                              mul_add[1][40]<=((mult_out_10[40] + mult_out_11[40] + mult_out_12[40])%3329) ;
                                                                              mul_add[1][41]<=((mult_out_10[41] + mult_out_11[41] + mult_out_12[41])%3329) ;
                                                                              mul_add[1][42]<=((mult_out_10[42] + mult_out_11[42] + mult_out_12[42])%3329) ;
                                                                              mul_add[1][43]<=((mult_out_10[43] + mult_out_11[43] + mult_out_12[43])%3329) ;
                                                                              mul_add[1][44]<=((mult_out_10[44] + mult_out_11[44] + mult_out_12[44])%3329) ;
                                                                              mul_add[1][45]<=((mult_out_10[45] + mult_out_11[45] + mult_out_12[45])%3329) ;
                                                                              mul_add[1][46]<=((mult_out_10[46] + mult_out_11[46] + mult_out_12[46])%3329) ;
                                                                              mul_add[1][47]<=((mult_out_10[47] + mult_out_11[47] + mult_out_12[47])%3329) ;
                                                                              mul_add[1][48]<=((mult_out_10[48] + mult_out_11[48] + mult_out_12[48])%3329) ;
                                                                              mul_add[1][49]<=((mult_out_10[49] + mult_out_11[49] + mult_out_12[49])%3329) ;
                                                                              mul_add[1][50]<=((mult_out_10[50] + mult_out_11[50] + mult_out_12[50])%3329) ;
                                                                              mul_add[1][51]<=((mult_out_10[51] + mult_out_11[51] + mult_out_12[51])%3329) ;
                                                                              mul_add[1][52]<=((mult_out_10[52] + mult_out_11[52] + mult_out_12[52])%3329) ;
                                                                              mul_add[1][53]<=((mult_out_10[53] + mult_out_11[53] + mult_out_12[53])%3329) ;
                                                                              mul_add[1][54]<=((mult_out_10[54] + mult_out_11[54] + mult_out_12[54])%3329) ;
                                                                              mul_add[1][55]<=((mult_out_10[55] + mult_out_11[55] + mult_out_12[55])%3329) ;
                                                                              mul_add[1][56]<=((mult_out_10[56] + mult_out_11[56] + mult_out_12[56])%3329) ;
                                                                              mul_add[1][57]<=((mult_out_10[57] + mult_out_11[57] + mult_out_12[57])%3329) ;
                                                                              mul_add[1][58]<=((mult_out_10[58] + mult_out_11[58] + mult_out_12[58])%3329) ;
                                                                              mul_add[1][59]<=((mult_out_10[59] + mult_out_11[59] + mult_out_12[59])%3329) ;
                                                                              mul_add[1][60]<=((mult_out_10[60] + mult_out_11[60] + mult_out_12[60])%3329) ;
                                                                              mul_add[1][61]<=((mult_out_10[61] + mult_out_11[61] + mult_out_12[61])%3329) ;
                                                                              mul_add[1][62]<=((mult_out_10[62] + mult_out_11[62] + mult_out_12[62])%3329) ;
                                                                              mul_add[1][63]<=((mult_out_10[63] + mult_out_11[63] + mult_out_12[63])%3329) ;
                                                                              mul_add[1][64]<=((mult_out_10[64] + mult_out_11[64] + mult_out_12[64])%3329) ;
                                                                              mul_add[1][65]<=((mult_out_10[65] + mult_out_11[65] + mult_out_12[65])%3329) ;
                                                                              mul_add[1][66]<=((mult_out_10[66] + mult_out_11[66] + mult_out_12[66])%3329) ;
                                                                              mul_add[1][67]<=((mult_out_10[67] + mult_out_11[67] + mult_out_12[67])%3329) ;
                                                                              mul_add[1][68]<=((mult_out_10[68] + mult_out_11[68] + mult_out_12[68])%3329) ;
                                                                              mul_add[1][69]<=((mult_out_10[69] + mult_out_11[69] + mult_out_12[69])%3329) ;
                                                                              mul_add[1][70]<=((mult_out_10[70] + mult_out_11[70] + mult_out_12[70])%3329) ;
                                                                              mul_add[1][71]<=((mult_out_10[71] + mult_out_11[71] + mult_out_12[71])%3329) ;
                                                                              mul_add[1][72]<=((mult_out_10[72] + mult_out_11[72] + mult_out_12[72])%3329) ;
                                                                              mul_add[1][73]<=((mult_out_10[73] + mult_out_11[73] + mult_out_12[73])%3329) ;
                                                                              mul_add[1][74]<=((mult_out_10[74] + mult_out_11[74] + mult_out_12[74])%3329) ;
                                                                              mul_add[1][75]<=((mult_out_10[75] + mult_out_11[75] + mult_out_12[75])%3329) ;
                                                                              mul_add[1][76]<=((mult_out_10[76] + mult_out_11[76] + mult_out_12[76])%3329) ;
                                                                              mul_add[1][77]<=((mult_out_10[77] + mult_out_11[77] + mult_out_12[77])%3329) ;
                                                                              mul_add[1][78]<=((mult_out_10[78] + mult_out_11[78] + mult_out_12[78])%3329) ;
                                                                              mul_add[1][79]<=((mult_out_10[79] + mult_out_11[79] + mult_out_12[79])%3329) ;
                                                                              mul_add[1][80]<=((mult_out_10[80] + mult_out_11[80] + mult_out_12[80])%3329) ;
                                                                              mul_add[1][81]<=((mult_out_10[81] + mult_out_11[81] + mult_out_12[81])%3329) ;
                                                                              mul_add[1][82]<=((mult_out_10[82] + mult_out_11[82] + mult_out_12[82])%3329) ;
                                                                              mul_add[1][83]<=((mult_out_10[83] + mult_out_11[83] + mult_out_12[83])%3329) ;
                                                                              mul_add[1][84]<=((mult_out_10[84] + mult_out_11[84] + mult_out_12[84])%3329) ;
                                                                              mul_add[1][85]<=((mult_out_10[85] + mult_out_11[85] + mult_out_12[85])%3329) ;
                                                                              mul_add[1][86]<=((mult_out_10[86] + mult_out_11[86] + mult_out_12[86])%3329) ;
                                                                              mul_add[1][87]<=((mult_out_10[87] + mult_out_11[87] + mult_out_12[87])%3329) ;
                                                                              mul_add[1][88]<=((mult_out_10[88] + mult_out_11[88] + mult_out_12[88])%3329) ;
                                                                              mul_add[1][89]<=((mult_out_10[89] + mult_out_11[89] + mult_out_12[89])%3329) ;
                                                                              mul_add[1][90]<=((mult_out_10[90] + mult_out_11[90] + mult_out_12[90])%3329) ;
                                                                              mul_add[1][91]<=((mult_out_10[91] + mult_out_11[91] + mult_out_12[91])%3329) ;
                                                                              mul_add[1][92]<=((mult_out_10[92] + mult_out_11[92] + mult_out_12[92])%3329) ;
                                                                              mul_add[1][93]<=((mult_out_10[93] + mult_out_11[93] + mult_out_12[93])%3329) ;
                                                                              mul_add[1][94]<=((mult_out_10[94] + mult_out_11[94] + mult_out_12[94])%3329) ;
                                                                              mul_add[1][95]<=((mult_out_10[95] + mult_out_11[95] + mult_out_12[95])%3329) ;
                                                                              mul_add[1][96]<=((mult_out_10[96] + mult_out_11[96] + mult_out_12[96])%3329) ;
                                                                              mul_add[1][97]<=((mult_out_10[97] + mult_out_11[97] + mult_out_12[97])%3329) ;
                                                                              mul_add[1][98]<=((mult_out_10[98] + mult_out_11[98] + mult_out_12[98])%3329) ;
                                                                              mul_add[1][99]<=((mult_out_10[99] + mult_out_11[99] + mult_out_12[99])%3329) ;
                                                                              mul_add[1][100]<=((mult_out_10[100] + mult_out_11[100] + mult_out_12[100])%3329);
                                                                              mul_add[1][101]<=((mult_out_10[101] + mult_out_11[101] + mult_out_12[101])%3329) ;
                                                                              mul_add[1][102]<=((mult_out_10[102] + mult_out_11[102] + mult_out_12[102])%3329) ;
                                                                              mul_add[1][103]<=((mult_out_10[103] + mult_out_11[103] + mult_out_12[103])%3329) ;
                                                                              mul_add[1][104]<=((mult_out_10[104] + mult_out_11[104] + mult_out_12[104])%3329) ;
                                                                              mul_add[1][105]<=((mult_out_10[105] + mult_out_11[105] + mult_out_12[105])%3329) ;
                                                                              mul_add[1][106]<=((mult_out_10[106] + mult_out_11[106] + mult_out_12[106])%3329) ;
                                                                              mul_add[1][107]<=((mult_out_10[107] + mult_out_11[107] + mult_out_12[107])%3329) ;
                                                                              mul_add[1][108]<=((mult_out_10[108] + mult_out_11[108] + mult_out_12[108])%3329) ;
                                                                              mul_add[1][109]<=((mult_out_10[109] + mult_out_11[109] + mult_out_12[109])%3329) ;
                                                                              mul_add[1][110]<=((mult_out_10[110] + mult_out_11[110] + mult_out_12[110])%3329) ;
                                                                              mul_add[1][111]<=((mult_out_10[111] + mult_out_11[111] + mult_out_12[111])%3329) ;
                                                                              mul_add[1][112]<=((mult_out_10[112] + mult_out_11[112] + mult_out_12[112])%3329) ;
                                                                              mul_add[1][113]<=((mult_out_10[113] + mult_out_11[113] + mult_out_12[113])%3329) ;
                                                                              mul_add[1][114]<=((mult_out_10[114] + mult_out_11[114] + mult_out_12[114])%3329) ;
                                                                              mul_add[1][115]<=((mult_out_10[115] + mult_out_11[115] + mult_out_12[115])%3329) ;
                                                                              mul_add[1][116]<=((mult_out_10[116] + mult_out_11[116] + mult_out_12[116])%3329) ;
                                                                              mul_add[1][117]<=((mult_out_10[117] + mult_out_11[117] + mult_out_12[117])%3329) ;
                                                                              mul_add[1][118]<=((mult_out_10[118] + mult_out_11[118] + mult_out_12[118])%3329) ;
                                                                              mul_add[1][119]<=((mult_out_10[119] + mult_out_11[119] + mult_out_12[119])%3329) ;
                                                                              mul_add[1][120]<=((mult_out_10[120] + mult_out_11[120] + mult_out_12[120])%3329) ;
                                                                              mul_add[1][121]<=((mult_out_10[121] + mult_out_11[121] + mult_out_12[121])%3329) ;
                                                                              mul_add[1][122]<=((mult_out_10[122] + mult_out_11[122] + mult_out_12[122])%3329) ;
                                                                              mul_add[1][123]<=((mult_out_10[123] + mult_out_11[123] + mult_out_12[123])%3329);
                                                                              mul_add[1][124]<=((mult_out_10[124] + mult_out_11[124] + mult_out_12[124])%3329);
                                                                              mul_add[1][125]<=((mult_out_10[125] + mult_out_11[125] + mult_out_12[125])%3329);
                                                                              mul_add[1][126]<=((mult_out_10[126] + mult_out_11[126] + mult_out_12[126])%3329);
                                                                              mul_add[1][127]<=((mult_out_10[127] + mult_out_11[127] + mult_out_12[127])%3329);
                                                                              mul_add[1][128]<=((mult_out_10[128] + mult_out_11[128] + mult_out_12[128])%3329);
                                                                              mul_add[1][129]<=((mult_out_10[129] + mult_out_11[129] + mult_out_12[129])%3329);
                                                                              mul_add[1][130]<=((mult_out_10[130] + mult_out_11[130] + mult_out_12[130])%3329);
                                                                              mul_add[1][131]<=((mult_out_10[131] + mult_out_11[131] + mult_out_12[131])%3329);
                                                                              mul_add[1][132]<=((mult_out_10[132] + mult_out_11[132] + mult_out_12[132])%3329);
                                                                              mul_add[1][133]<=((mult_out_10[133] + mult_out_11[133] + mult_out_12[133])%3329);
                                                                              mul_add[1][134]<=((mult_out_10[134] + mult_out_11[134] + mult_out_12[134])%3329);
                                                                              mul_add[1][135]<=((mult_out_10[135] + mult_out_11[135] + mult_out_12[135])%3329);
                                                                              mul_add[1][136]<=((mult_out_10[136] + mult_out_11[136] + mult_out_12[136])%3329);
                                                                              mul_add[1][137]<=((mult_out_10[137] + mult_out_11[137] + mult_out_12[137])%3329);
                                                                              mul_add[1][138]<=((mult_out_10[138] + mult_out_11[138] + mult_out_12[138])%3329);
                                                                              mul_add[1][139]<=((mult_out_10[139] + mult_out_11[139] + mult_out_12[139])%3329);
                                                                              mul_add[1][140]<=((mult_out_10[140] + mult_out_11[140] + mult_out_12[140])%3329);
                                                                              mul_add[1][141]<=((mult_out_10[141] + mult_out_11[141] + mult_out_12[141])%3329);
                                                                              mul_add[1][142]<=((mult_out_10[142] + mult_out_11[142] + mult_out_12[142])%3329);
                                                                              mul_add[1][143]<=((mult_out_10[143] + mult_out_11[143] + mult_out_12[143])%3329);
                                                                              mul_add[1][144]<=((mult_out_10[144] + mult_out_11[144] + mult_out_12[144])%3329);
                                                                              mul_add[1][145]<=((mult_out_10[145] + mult_out_11[145] + mult_out_12[145])%3329);
                                                                              mul_add[1][146]<=((mult_out_10[146] + mult_out_11[146] + mult_out_12[146])%3329);
                                                                              mul_add[1][147]<=((mult_out_10[147] + mult_out_11[147] + mult_out_12[147])%3329);
                                                                              mul_add[1][148]<=((mult_out_10[148] + mult_out_11[148] + mult_out_12[148])%3329);
                                                                              mul_add[1][149]<=((mult_out_10[149] + mult_out_11[149] + mult_out_12[149])%3329);
                                                                              mul_add[1][150]<=((mult_out_10[150] + mult_out_11[150] + mult_out_12[150])%3329);
                                                                              mul_add[1][151]<=((mult_out_10[151] + mult_out_11[151] + mult_out_12[151])%3329);
                                                                              mul_add[1][152]<=((mult_out_10[152] + mult_out_11[152] + mult_out_12[152])%3329);
                                                                              mul_add[1][153]<=((mult_out_10[153] + mult_out_11[153] + mult_out_12[153])%3329);
                                                                              mul_add[1][154]<=((mult_out_10[154] + mult_out_11[154] + mult_out_12[154])%3329);
                                                                              mul_add[1][155]<=((mult_out_10[155] + mult_out_11[155] + mult_out_12[155])%3329);
                                                                              mul_add[1][156]<=((mult_out_10[156] + mult_out_11[156] + mult_out_12[156])%3329);
                                                                              mul_add[1][157]<=((mult_out_10[157] + mult_out_11[157] + mult_out_12[157])%3329) ;
                                                                              mul_add[1][158]<=((mult_out_10[158] + mult_out_11[158] + mult_out_12[158])%3329) ;
                                                                              mul_add[1][159]<=((mult_out_10[159] + mult_out_11[159] + mult_out_12[159])%3329);
                                                                              mul_add[1][160]<=((mult_out_10[160] + mult_out_11[160] + mult_out_12[160])%3329) ;
                                                                              mul_add[1][161]<=((mult_out_10[161] + mult_out_11[161] + mult_out_12[161])%3329) ;
                                                                              mul_add[1][162]<=((mult_out_10[162] + mult_out_11[162] + mult_out_12[162])%3329) ;
                                                                              mul_add[1][163]<=((mult_out_10[163] + mult_out_11[163] + mult_out_12[163])%3329);
                                                                              mul_add[1][164]<=((mult_out_10[164] + mult_out_11[164] + mult_out_12[164])%3329);
                                                                              mul_add[1][165]<=((mult_out_10[165] + mult_out_11[165] + mult_out_12[165])%3329) ;
                                                                              mul_add[1][166]<=((mult_out_10[166] + mult_out_11[166] + mult_out_12[166])%3329) ;
                                                                              mul_add[1][167]<=((mult_out_10[167] + mult_out_11[167] + mult_out_12[167])%3329) ;
                                                                              mul_add[1][168]<=((mult_out_10[168] + mult_out_11[168] + mult_out_12[168])%3329) ;
                                                                              mul_add[1][169]<=((mult_out_10[169] + mult_out_11[169] + mult_out_12[169])%3329) ;
                                                                              mul_add[1][170]<=((mult_out_10[170] + mult_out_11[170] + mult_out_12[170])%3329) ;
                                                                              mul_add[1][171]<=((mult_out_10[171] + mult_out_11[171] + mult_out_12[171])%3329) ;
                                                                              mul_add[1][172]<=((mult_out_10[172] + mult_out_11[172] + mult_out_12[172])%3329) ;
                                                                              mul_add[1][173]<=((mult_out_10[173] + mult_out_11[173] + mult_out_12[173])%3329) ;
                                                                              mul_add[1][174]<=((mult_out_10[174] + mult_out_11[174] + mult_out_12[174])%3329) ;
                                                                              mul_add[1][175]<=((mult_out_10[175] + mult_out_11[175] + mult_out_12[175])%3329) ;
                                                                              mul_add[1][176]<=((mult_out_10[176] + mult_out_11[176] + mult_out_12[176])%3329) ;
                                                                              mul_add[1][177]<=((mult_out_10[177] + mult_out_11[177] + mult_out_12[177])%3329) ;
                                                                              mul_add[1][178]<=((mult_out_10[178] + mult_out_11[178] + mult_out_12[178])%3329) ;
                                                                              mul_add[1][179]<=((mult_out_10[179] + mult_out_11[179] + mult_out_12[179])%3329) ;
                                                                              mul_add[1][180]<=((mult_out_10[180] + mult_out_11[180] + mult_out_12[180])%3329) ;
                                                                              mul_add[1][181]<=((mult_out_10[181] + mult_out_11[181] + mult_out_12[181])%3329) ;
                                                                              mul_add[1][182]<=((mult_out_10[182] + mult_out_11[182] + mult_out_12[182])%3329) ;
                                                                              mul_add[1][183]<=((mult_out_10[183] + mult_out_11[183] + mult_out_12[183])%3329) ;
                                                                              mul_add[1][184]<=((mult_out_10[184] + mult_out_11[184] + mult_out_12[184])%3329) ;
                                                                              mul_add[1][185]<=((mult_out_10[185] + mult_out_11[185] + mult_out_12[185])%3329) ;
                                                                              mul_add[1][186]<=((mult_out_10[186] + mult_out_11[186] + mult_out_12[186])%3329) ;
                                                                              mul_add[1][187]<=((mult_out_10[187] + mult_out_11[187] + mult_out_12[187])%3329) ;
                                                                              mul_add[1][188]<=((mult_out_10[188] + mult_out_11[188] + mult_out_12[188])%3329) ;
                                                                              mul_add[1][189]<=((mult_out_10[189] + mult_out_11[189] + mult_out_12[189])%3329) ;
                                                                              mul_add[1][190]<=((mult_out_10[190] + mult_out_11[190] + mult_out_12[190])%3329) ;
                                                                              mul_add[1][191]<=((mult_out_10[191] + mult_out_11[191] + mult_out_12[191])%3329) ;
                                                                              mul_add[1][192]<=((mult_out_10[192] + mult_out_11[192] + mult_out_12[192])%3329) ;
                                                                              mul_add[1][193]<=((mult_out_10[193] + mult_out_11[193] + mult_out_12[193])%3329) ;
                                                                              mul_add[1][194]<=((mult_out_10[194] + mult_out_11[194] + mult_out_12[194])%3329) ;
                                                                              mul_add[1][195]<=((mult_out_10[195] + mult_out_11[195] + mult_out_12[195])%3329) ;
                                                                              mul_add[1][196]<=((mult_out_10[196] + mult_out_11[196] + mult_out_12[196])%3329) ;
                                                                              mul_add[1][197]<=((mult_out_10[197] + mult_out_11[197] + mult_out_12[197])%3329) ;
                                                                              mul_add[1][198]<=((mult_out_10[198] + mult_out_11[198] + mult_out_12[198])%3329) ;
                                                                              mul_add[1][199]<=((mult_out_10[199] + mult_out_11[199] + mult_out_12[199])%3329) ;
                                                                              mul_add[1][200]<=((mult_out_10[200] + mult_out_11[200] + mult_out_12[200])%3329) ;
                                                                              mul_add[1][201]<=((mult_out_10[201] + mult_out_11[201] + mult_out_12[201])%3329) ;
                                                                              mul_add[1][202]<=((mult_out_10[202] + mult_out_11[202] + mult_out_12[202])%3329) ;
                                                                              mul_add[1][203]<=((mult_out_10[203] + mult_out_11[203] + mult_out_12[203])%3329) ;
                                                                              mul_add[1][204]<=((mult_out_10[204] + mult_out_11[204] + mult_out_12[204])%3329) ;
                                                                              mul_add[1][205]<=((mult_out_10[205] + mult_out_11[205] + mult_out_12[205])%3329) ;
                                                                              mul_add[1][206]<=((mult_out_10[206] + mult_out_11[206] + mult_out_12[206])%3329) ;
                                                                              mul_add[1][207]<=((mult_out_10[207] + mult_out_11[207] + mult_out_12[207])%3329) ;
                                                                              mul_add[1][208]<=((mult_out_10[208] + mult_out_11[208] + mult_out_12[208])%3329) ;
                                                                              mul_add[1][209]<=((mult_out_10[209] + mult_out_11[209] + mult_out_12[209])%3329) ;
                                                                              mul_add[1][210]<=((mult_out_10[210] + mult_out_11[210] + mult_out_12[210])%3329) ;
                                                                              mul_add[1][211]<=((mult_out_10[211] + mult_out_11[211] + mult_out_12[211])%3329) ;
                                                                              mul_add[1][212]<=((mult_out_10[212] + mult_out_11[212] + mult_out_12[212])%3329) ;
                                                                              mul_add[1][213]<=((mult_out_10[213] + mult_out_11[213] + mult_out_12[213])%3329) ;
                                                                              mul_add[1][214]<=((mult_out_10[214] + mult_out_11[214] + mult_out_12[214])%3329) ;
                                                                              mul_add[1][215]<=((mult_out_10[215] + mult_out_11[215] + mult_out_12[215])%3329) ;
                                                                              mul_add[1][216]<=((mult_out_10[216] + mult_out_11[216] + mult_out_12[216])%3329) ;
                                                                              mul_add[1][217]<=((mult_out_10[217] + mult_out_11[217] + mult_out_12[217])%3329) ;
                                                                              mul_add[1][218]<=((mult_out_10[218] + mult_out_11[218] + mult_out_12[218])%3329) ;
                                                                              mul_add[1][219]<=((mult_out_10[219] + mult_out_11[219] + mult_out_12[219])%3329) ;
                                                                              mul_add[1][220]<=((mult_out_10[220] + mult_out_11[220] + mult_out_12[220])%3329) ;
                                                                              mul_add[1][221]<=((mult_out_10[221] + mult_out_11[221] + mult_out_12[221])%3329) ;
                                                                              mul_add[1][222]<=((mult_out_10[222] + mult_out_11[222] + mult_out_12[222])%3329) ;
                                                                              mul_add[1][223]<=((mult_out_10[223] + mult_out_11[223] + mult_out_12[223])%3329) ;
                                                                              mul_add[1][224]<=((mult_out_10[224] + mult_out_11[224] + mult_out_12[224])%3329) ;
                                                                              mul_add[1][225]<=((mult_out_10[225] + mult_out_11[225] + mult_out_12[225])%3329) ;
                                                                              mul_add[1][226]<=((mult_out_10[226] + mult_out_11[226] + mult_out_12[226])%3329) ;
                                                                              mul_add[1][227]<=((mult_out_10[227] + mult_out_11[227] + mult_out_12[227])%3329) ;
                                                                              mul_add[1][228]<=((mult_out_10[228] + mult_out_11[228] + mult_out_12[228])%3329) ;
                                                                              mul_add[1][229]<=((mult_out_10[229] + mult_out_11[229] + mult_out_12[229])%3329) ;
                                                                              mul_add[1][230]<=((mult_out_10[230] + mult_out_11[230] + mult_out_12[230])%3329) ;
                                                                              mul_add[1][231]<=((mult_out_10[231] + mult_out_11[231] + mult_out_12[231])%3329) ;
                                                                              mul_add[1][232]<=((mult_out_10[232] + mult_out_11[232] + mult_out_12[232])%3329) ;
                                                                              mul_add[1][233]<=((mult_out_10[233] + mult_out_11[233] + mult_out_12[233])%3329) ;
                                                                              mul_add[1][234]<=((mult_out_10[234] + mult_out_11[234] + mult_out_12[234])%3329) ;
                                                                              mul_add[1][235]<=((mult_out_10[235] + mult_out_11[235] + mult_out_12[235])%3329) ;
                                                                              mul_add[1][236]<=((mult_out_10[236] + mult_out_11[236] + mult_out_12[236])%3329) ;
                                                                              mul_add[1][237]<=((mult_out_10[237] + mult_out_11[237] + mult_out_12[237])%3329) ;
                                                                              mul_add[1][238]<=((mult_out_10[238] + mult_out_11[238] + mult_out_12[238])%3329) ;
                                                                              mul_add[1][239]<=((mult_out_10[239] + mult_out_11[239] + mult_out_12[239])%3329) ;
                                                                              mul_add[1][240]<=((mult_out_10[240] + mult_out_11[240] + mult_out_12[240])%3329) ;
                                                                              mul_add[1][241]<=((mult_out_10[241] + mult_out_11[241] + mult_out_12[241])%3329) ;
                                                                              mul_add[1][242]<=((mult_out_10[242] + mult_out_11[242] + mult_out_12[242])%3329) ;
                                                                              mul_add[1][243]<=((mult_out_10[243] + mult_out_11[243] + mult_out_12[243])%3329) ;
                                                                              mul_add[1][244]<=((mult_out_10[244] + mult_out_11[244] + mult_out_12[244])%3329) 
                                                                              mul_add[1][245]<=((mult_out_10[245] + mult_out_11[245] + mult_out_12[245])%3329) ;
                                                                              mul_add[1][246]<=((mult_out_10[246] + mult_out_11[246] + mult_out_12[246])%3329) ;
                                                                              mul_add[1][247]<=((mult_out_10[247] + mult_out_11[247] + mult_out_12[247])%3329);
                                                                              mul_add[1][248]<=((mult_out_10[248] + mult_out_11[248] + mult_out_12[248])%3329) ;
                                                                              mul_add[1][249]<=((mult_out_10[249] + mult_out_11[249] + mult_out_12[249])%3329) ;
                                                                              mul_add[1][250]<=((mult_out_10[250] + mult_out_11[250] + mult_out_12[250])%3329) ;
                                                                              mul_add[1][251]<=((mult_out_10[251] + mult_out_11[251] + mult_out_12[251])%3329) ;
                                                                              mul_add[1][252]<=((mult_out_10[252] + mult_out_11[252] + mult_out_12[252])%3329) ;
                                                                              mul_add[1][253]<=((mult_out_10[253] + mult_out_11[253] + mult_out_12[253])%3329) ;
                                                                              mul_add[1][254]<=((mult_out_10[254] + mult_out_11[254] + mult_out_12[254])%3329) ;
                                                                              mul_add[1][255]<=((mult_out_10[255] + mult_out_11[255] + mult_out_12[255])%3329) ;
                                                                             
                                                                         
                                                                              mul_add[2][0]<=((mult_out_20[0] + mult_out_21[0] + mult_out_22[0])%3329) ;
                                                                          mul_add[2][1]<=((mult_out_20[1] + mult_out_21[1] + mult_out_22[1])%3329) ;
                                                                          mul_add[2][2]<=((mult_out_20[2] + mult_out_21[2] + mult_out_22[2])%3329) ;
                                                                          mul_add[2][3]<=((mult_out_20[3] + mult_out_21[3] + mult_out_22[3])%3329) ;
                                                                          mul_add[2][4]<=((mult_out_20[4] + mult_out_21[4] + mult_out_22[4])%3329) ;
                                                                          mul_add[2][5]<=((mult_out_20[5] + mult_out_21[5] + mult_out_22[5])%3329) ;
                                                                          mul_add[2][6]<=((mult_out_20[6] + mult_out_21[6] + mult_out_22[6])%3329) ;
                                                                          mul_add[2][7]<=((mult_out_20[7] + mult_out_21[7] + mult_out_22[7])%3329) ;
                                                                          mul_add[2][8]<=((mult_out_20[8] + mult_out_21[8] + mult_out_22[8])%3329) ;
                                                                          mul_add[2][9]<=((mult_out_20[9] + mult_out_21[9] + mult_out_22[9])%3329) ;
                                                                          mul_add[2][10]<=((mult_out_20[10] + mult_out_21[10] + mult_out_22[10])%3329) ;
                                                                          mul_add[2][11]<=((mult_out_20[11] + mult_out_21[11] + mult_out_22[11])%3329) ;
                                                                          mul_add[2][12]<=((mult_out_20[12] + mult_out_21[12] + mult_out_22[12])%3329) ;
                                                                          mul_add[2][13]<=((mult_out_20[13] + mult_out_21[13] + mult_out_22[13])%3329) ;
                                                                          mul_add[2][14]<=((mult_out_20[14] + mult_out_21[14] + mult_out_22[14])%3329) ;
                                                                          mul_add[2][15]<=((mult_out_20[15] + mult_out_21[15] + mult_out_22[15])%3329) ;
                                                                          mul_add[2][16]<=((mult_out_20[16] + mult_out_21[16] + mult_out_22[16])%3329) ;
                                                                          mul_add[2][17]<=((mult_out_20[17] + mult_out_21[17] + mult_out_22[17])%3329) ;
                                                                          mul_add[2][18]<=((mult_out_20[18] + mult_out_21[18] + mult_out_22[18])%3329) ;
                                                                          mul_add[2][19]<=((mult_out_20[19] + mult_out_21[19] + mult_out_22[19])%3329) ;
                                                                          mul_add[2][20]<=((mult_out_20[20] + mult_out_21[20] + mult_out_22[20])%3329) ;
                                                                          mul_add[2][21]<=((mult_out_20[21] + mult_out_21[21] + mult_out_22[21])%3329) ;
                                                                          mul_add[2][22]<=((mult_out_20[22] + mult_out_21[22] + mult_out_22[22])%3329) ;
                                                                          mul_add[2][23]<=((mult_out_20[23] + mult_out_21[23] + mult_out_22[23])%3329) ;
                                                                          mul_add[2][24]<=((mult_out_20[24] + mult_out_21[24] + mult_out_22[24])%3329) ;
                                                                          mul_add[2][25]<=((mult_out_20[25] + mult_out_21[25] + mult_out_22[25])%3329) ;
                                                                          mul_add[2][26]<=((mult_out_20[26] + mult_out_21[26] + mult_out_22[26])%3329) ;
                                                                          mul_add[2][27]<=((mult_out_20[27] + mult_out_21[27] + mult_out_22[27])%3329) ;
                                                                          mul_add[2][28]<=((mult_out_20[28] + mult_out_21[28] + mult_out_22[28])%3329) ;
                                                                          mul_add[2][29]<=((mult_out_20[29] + mult_out_21[29] + mult_out_22[29])%3329) ;
                                                                          mul_add[2][30]<=((mult_out_20[30] + mult_out_21[30] + mult_out_22[30])%3329) ;
                                                                          mul_add[2][31]<=((mult_out_20[31] + mult_out_21[31] + mult_out_22[31])%3329) ;
                                                                          mul_add[2][32]<=((mult_out_20[32] + mult_out_21[32] + mult_out_22[32])%3329) ;
                                                                          mul_add[2][33]<=((mult_out_20[33] + mult_out_21[33] + mult_out_22[33])%3329) ;
                                                                          mul_add[2][34]<=((mult_out_20[34] + mult_out_21[34] + mult_out_22[34])%3329) ;
                                                                          mul_add[2][35]<=((mult_out_20[35] + mult_out_21[35] + mult_out_22[35])%3329) ;
                                                                          mul_add[2][36]<=((mult_out_20[36] + mult_out_21[36] + mult_out_22[36])%3329) ;
                                                                          mul_add[2][37]<=((mult_out_20[37] + mult_out_21[37] + mult_out_22[37])%3329) ;
                                                                          mul_add[2][38]<=((mult_out_20[38] + mult_out_21[38] + mult_out_22[38])%3329) ;
                                                                          mul_add[2][39]<=((mult_out_20[39] + mult_out_21[39] + mult_out_22[39])%3329) ;
                                                                          mul_add[2][40]<=((mult_out_20[40] + mult_out_21[40] + mult_out_22[40])%3329) ;
                                                                          mul_add[2][41]<=((mult_out_20[41] + mult_out_21[41] + mult_out_22[41])%3329) ;
                                                                          mul_add[2][42]<=((mult_out_20[42] + mult_out_21[42] + mult_out_22[42])%3329) ;
                                                                          mul_add[2][43]<=((mult_out_20[43] + mult_out_21[43] + mult_out_22[43])%3329) ;
                                                                          mul_add[2][44]<=((mult_out_20[44] + mult_out_21[44] + mult_out_22[44])%3329) ;
                                                                          mul_add[2][45]<=((mult_out_20[45] + mult_out_21[45] + mult_out_22[45])%3329) ;
                                                                          mul_add[2][46]<=((mult_out_20[46] + mult_out_21[46] + mult_out_22[46])%3329) ;
                                                                          mul_add[2][47]<=((mult_out_20[47] + mult_out_21[47] + mult_out_22[47])%3329) ;
                                                                          mul_add[2][48]<=((mult_out_20[48] + mult_out_21[48] + mult_out_22[48])%3329) ;
                                                                          mul_add[2][49]<=((mult_out_20[49] + mult_out_21[49] + mult_out_22[49])%3329) ;
                                                                          mul_add[2][50]<=((mult_out_20[50] + mult_out_21[50] + mult_out_22[50])%3329) ;
                                                                          mul_add[2][51]<=((mult_out_20[51] + mult_out_21[51] + mult_out_22[51])%3329) ;
                                                                          mul_add[2][52]<=((mult_out_20[52] + mult_out_21[52] + mult_out_22[52])%3329) ;
                                                                          mul_add[2][53]<=((mult_out_20[53] + mult_out_21[53] + mult_out_22[53])%3329) ;
                                                                          mul_add[2][54]<=((mult_out_20[54] + mult_out_21[54] + mult_out_22[54])%3329) ;
                                                                          mul_add[2][55]<=((mult_out_20[55] + mult_out_21[55] + mult_out_22[55])%3329) ;
                                                                          mul_add[2][56]<=((mult_out_20[56] + mult_out_21[56] + mult_out_22[56])%3329) ;
                                                                          mul_add[2][57]<=((mult_out_20[57] + mult_out_21[57] + mult_out_22[57])%3329) ;
                                                                          mul_add[2][58]<=((mult_out_20[58] + mult_out_21[58] + mult_out_22[58])%3329) ;
                                                                          mul_add[2][59]<=((mult_out_20[59] + mult_out_21[59] + mult_out_22[59])%3329) ;
                                                                          mul_add[2][60]<=((mult_out_20[60] + mult_out_21[60] + mult_out_22[60])%3329) ;
                                                                          mul_add[2][61]<=((mult_out_20[61] + mult_out_21[61] + mult_out_22[61])%3329) ;
                                                                          mul_add[2][62]<=((mult_out_20[62] + mult_out_21[62] + mult_out_22[62])%3329) ;
                                                                          mul_add[2][63]<=((mult_out_20[63] + mult_out_21[63] + mult_out_22[63])%3329) ;
                                                                          mul_add[2][64]<=((mult_out_20[64] + mult_out_21[64] + mult_out_22[64])%3329) ;
                                                                          mul_add[2][65]<=((mult_out_20[65] + mult_out_21[65] + mult_out_22[65])%3329) ;
                                                                          mul_add[2][66]<=((mult_out_20[66] + mult_out_21[66] + mult_out_22[66])%3329) ;
                                                                          mul_add[2][67]<=((mult_out_20[67] + mult_out_21[67] + mult_out_22[67])%3329) ;
                                                                          mul_add[2][68]<=((mult_out_20[68] + mult_out_21[68] + mult_out_22[68])%3329) ;
                                                                          mul_add[2][69]<=((mult_out_20[69] + mult_out_21[69] + mult_out_22[69])%3329) ;
                                                                          mul_add[2][70]<=((mult_out_20[70] + mult_out_21[70] + mult_out_22[70])%3329) ;
                                                                          mul_add[2][71]<=((mult_out_20[71] + mult_out_21[71] + mult_out_22[71])%3329) ;
                                                                          mul_add[2][72]<=((mult_out_20[72] + mult_out_21[72] + mult_out_22[72])%3329) ;
                                                                          mul_add[2][73]<=((mult_out_20[73] + mult_out_21[73] + mult_out_22[73])%3329) ;
                                                                          mul_add[2][74]<=((mult_out_20[74] + mult_out_21[74] + mult_out_22[74])%3329) ;
                                                                          mul_add[2][75]<=((mult_out_20[75] + mult_out_21[75] + mult_out_22[75])%3329) ;
                                                                          mul_add[2][76]<=((mult_out_20[76] + mult_out_21[76] + mult_out_22[76])%3329) ;
                                                                          mul_add[2][77]<=((mult_out_20[77] + mult_out_21[77] + mult_out_22[77])%3329) ;
                                                                          mul_add[2][78]<=((mult_out_20[78] + mult_out_21[78] + mult_out_22[78])%3329) ;
                                                                          mul_add[2][79]<=((mult_out_20[79] + mult_out_21[79] + mult_out_22[79])%3329) ;
                                                                          mul_add[2][80]<=((mult_out_20[80] + mult_out_21[80] + mult_out_22[80])%3329) ;
                                                                          mul_add[2][81]<=((mult_out_20[81] + mult_out_21[81] + mult_out_22[81])%3329) ;
                                                                          mul_add[2][82]<=((mult_out_20[82] + mult_out_21[82] + mult_out_22[82])%3329) ;
                                                                          mul_add[2][83]<=((mult_out_20[83] + mult_out_21[83] + mult_out_22[83])%3329) ;
                                                                          mul_add[2][84]<=((mult_out_20[84] + mult_out_21[84] + mult_out_22[84])%3329) ;
                                                                          mul_add[2][85]<=((mult_out_20[85] + mult_out_21[85] + mult_out_22[85])%3329) ;
                                                                          mul_add[2][86]<=((mult_out_20[86] + mult_out_21[86] + mult_out_22[86])%3329) ;
                                                                          mul_add[2][87]<=((mult_out_20[87] + mult_out_21[87] + mult_out_22[87])%3329) ;
                                                                          mul_add[2][88]<=((mult_out_20[88] + mult_out_21[88] + mult_out_22[88])%3329) ;
                                                                          mul_add[2][89]<=((mult_out_20[89] + mult_out_21[89] + mult_out_22[89])%3329) ;
                                                                          mul_add[2][90]<=((mult_out_20[90] + mult_out_21[90] + mult_out_22[90])%3329) ;
                                                                          mul_add[2][91]<=((mult_out_20[91] + mult_out_21[91] + mult_out_22[91])%3329) ;
                                                                          mul_add[2][92]<=((mult_out_20[92] + mult_out_21[92] + mult_out_22[92])%3329) ;
                                                                          mul_add[2][93]<=((mult_out_20[93] + mult_out_21[93] + mult_out_22[93])%3329) ;
                                                                          mul_add[2][94]<=((mult_out_20[94] + mult_out_21[94] + mult_out_22[94])%3329) ;
                                                                          mul_add[2][95]<=((mult_out_20[95] + mult_out_21[95] + mult_out_22[95])%3329) ;
                                                                          mul_add[2][96]<=((mult_out_20[96] + mult_out_21[96] + mult_out_22[96])%3329) ;
                                                                          mul_add[2][97]<=((mult_out_20[97] + mult_out_21[97] + mult_out_22[97])%3329) ;
                                                                          mul_add[2][98]<=((mult_out_20[98] + mult_out_21[98] + mult_out_22[98])%3329) ;
                                                                          mul_add[2][99]<=((mult_out_20[99] + mult_out_21[99] + mult_out_22[99])%3329) ;
                                                                          mul_add[2][100]<=((mult_out_20[100] + mult_out_21[100] + mult_out_22[100])%3329) ;
                                                                          mul_add[2][101]<=((mult_out_20[101] + mult_out_21[101] + mult_out_22[101])%3329) ;
                                                                          mul_add[2][102]<=((mult_out_20[102] + mult_out_21[102] + mult_out_22[102])%3329) ;
                                                                          mul_add[2][103]<=((mult_out_20[103] + mult_out_21[103] + mult_out_22[103])%3329) ;
                                                                          mul_add[2][104]<=((mult_out_20[104] + mult_out_21[104] + mult_out_22[104])%3329) ;
                                                                          mul_add[2][105]<=((mult_out_20[105] + mult_out_21[105] + mult_out_22[105])%3329) ;
                                                                          mul_add[2][106]<=((mult_out_20[106] + mult_out_21[106] + mult_out_22[106])%3329) ;
                                                                          mul_add[2][107]<=((mult_out_20[107] + mult_out_21[107] + mult_out_22[107])%3329) ;
                                                                          mul_add[2][108]<=((mult_out_20[108] + mult_out_21[108] + mult_out_22[108])%3329) ;
                                                                          mul_add[2][109]<=((mult_out_20[109] + mult_out_21[109] + mult_out_22[109])%3329) ;
                                                                          mul_add[2][110]<=((mult_out_20[110] + mult_out_21[110] + mult_out_22[110])%3329) ;
                                                                          mul_add[2][111]<=((mult_out_20[111] + mult_out_21[111] + mult_out_22[111])%3329) ;
                                                                          mul_add[2][112]<=((mult_out_20[112] + mult_out_21[112] + mult_out_22[112])%3329) ;
                                                                          mul_add[2][113]<=((mult_out_20[113] + mult_out_21[113] + mult_out_22[113])%3329) ;
                                                                          mul_add[2][114]<=((mult_out_20[114] + mult_out_21[114] + mult_out_22[114])%3329) ;
                                                                          mul_add[2][115]<=((mult_out_20[115] + mult_out_21[115] + mult_out_22[115])%3329) ;
                                                                          mul_add[2][116]<=((mult_out_20[116] + mult_out_21[116] + mult_out_22[116])%3329) ;
                                                                          mul_add[2][117]<=((mult_out_20[117] + mult_out_21[117] + mult_out_22[117])%3329) ;
                                                                          mul_add[2][118]<=((mult_out_20[118] + mult_out_21[118] + mult_out_22[118])%3329) ;
                                                                          mul_add[2][119]<=((mult_out_20[119] + mult_out_21[119] + mult_out_22[119])%3329) ;
                                                                          mul_add[2][120]<=((mult_out_20[120] + mult_out_21[120] + mult_out_22[120])%3329) ;
                                                                          mul_add[2][121]<=((mult_out_20[121] + mult_out_21[121] + mult_out_22[121])%3329) ;
                                                                          mul_add[2][122]<=((mult_out_20[122] + mult_out_21[122] + mult_out_22[122])%3329) ;
                                                                          mul_add[2][123]<=((mult_out_20[123] + mult_out_21[123] + mult_out_22[123])%3329) ;
                                                                          mul_add[2][124]<=((mult_out_20[124] + mult_out_21[124] + mult_out_22[124])%3329) ;
                                                                          mul_add[2][125]<=((mult_out_20[125] + mult_out_21[125] + mult_out_22[125])%3329) ;
                                                                          mul_add[2][126]<=((mult_out_20[126] + mult_out_21[126] + mult_out_22[126])%3329) ;
                                                                          mul_add[2][127]<=((mult_out_20[127] + mult_out_21[127] + mult_out_22[127])%3329) ;
                                                                          mul_add[2][128]<=((mult_out_20[128] + mult_out_21[128] + mult_out_22[128])%3329) ;
                                                                          mul_add[2][129]<=((mult_out_20[129] + mult_out_21[129] + mult_out_22[129])%3329) ;
                                                                          mul_add[2][130]<=((mult_out_20[130] + mult_out_21[130] + mult_out_22[130])%3329) ;
                                                                          mul_add[2][131]<=((mult_out_20[131] + mult_out_21[131] + mult_out_22[131])%3329) ;
                                                                          mul_add[2][132]<=((mult_out_20[132] + mult_out_21[132] + mult_out_22[132])%3329) ;
                                                                          mul_add[2][133]<=((mult_out_20[133] + mult_out_21[133] + mult_out_22[133])%3329) ;
                                                                          mul_add[2][134]<=((mult_out_20[134] + mult_out_21[134] + mult_out_22[134])%3329) ;
                                                                          mul_add[2][135]<=((mult_out_20[135] + mult_out_21[135] + mult_out_22[135])%3329) ;
                                                                          mul_add[2][136]<=((mult_out_20[136] + mult_out_21[136] + mult_out_22[136])%3329) ;
                                                                          mul_add[2][137]<=((mult_out_20[137] + mult_out_21[137] + mult_out_22[137])%3329) ;
                                                                          mul_add[2][138]<=((mult_out_20[138] + mult_out_21[138] + mult_out_22[138])%3329) ;
                                                                          mul_add[2][139]<=((mult_out_20[139] + mult_out_21[139] + mult_out_22[139])%3329) ;
                                                                          mul_add[2][140]<=((mult_out_20[140] + mult_out_21[140] + mult_out_22[140])%3329) ;
                                                                          mul_add[2][141]<=((mult_out_20[141] + mult_out_21[141] + mult_out_22[141])%3329) ;
                                                                          mul_add[2][142]<=((mult_out_20[142] + mult_out_21[142] + mult_out_22[142])%3329) ;
                                                                          mul_add[2][143]<=((mult_out_20[143] + mult_out_21[143] + mult_out_22[143])%3329) ;
                                                                          mul_add[2][144]<=((mult_out_20[144] + mult_out_21[144] + mult_out_22[144])%3329) ;
                                                                          mul_add[2][145]<=((mult_out_20[145] + mult_out_21[145] + mult_out_22[145])%3329) ;
                                                                          mul_add[2][146]<=((mult_out_20[146] + mult_out_21[146] + mult_out_22[146])%3329) ;
                                                                          mul_add[2][147]<=((mult_out_20[147] + mult_out_21[147] + mult_out_22[147])%3329) ;
                                                                          mul_add[2][148]<=((mult_out_20[148] + mult_out_21[148] + mult_out_22[148])%3329) ;
                                                                          mul_add[2][149]<=((mult_out_20[149] + mult_out_21[149] + mult_out_22[149])%3329) ;
                                                                          mul_add[2][150]<=((mult_out_20[150] + mult_out_21[150] + mult_out_22[150])%3329) ;
                                                                          mul_add[2][151]<=((mult_out_20[151] + mult_out_21[151] + mult_out_22[151])%3329) ;
                                                                          mul_add[2][152]<=((mult_out_20[152] + mult_out_21[152] + mult_out_22[152])%3329) ;
                                                                          mul_add[2][153]<=((mult_out_20[153] + mult_out_21[153] + mult_out_22[153])%3329) ;
                                                                          mul_add[2][154]<=((mult_out_20[154] + mult_out_21[154] + mult_out_22[154])%3329) ;
                                                                          mul_add[2][155]<=((mult_out_20[155] + mult_out_21[155] + mult_out_22[155])%3329) ;
                                                                          mul_add[2][156]<=((mult_out_20[156] + mult_out_21[156] + mult_out_22[156])%3329) ;
                                                                          mul_add[2][157]<=((mult_out_20[157] + mult_out_21[157] + mult_out_22[157])%3329) ;
                                                                          mul_add[2][158]<=((mult_out_20[158] + mult_out_21[158] + mult_out_22[158])%3329) ;
                                                                          mul_add[2][159]<=((mult_out_20[159] + mult_out_21[159] + mult_out_22[159])%3329) ;
                                                                          mul_add[2][160]<=((mult_out_20[160] + mult_out_21[160] + mult_out_22[160])%3329) ;
                                                                          mul_add[2][161]<=((mult_out_20[161] + mult_out_21[161] + mult_out_22[161])%3329) ;
                                                                          mul_add[2][162]<=((mult_out_20[162] + mult_out_21[162] + mult_out_22[162])%3329) ;
                                                                          mul_add[2][163]<=((mult_out_20[163] + mult_out_21[163] + mult_out_22[163])%3329) ;
                                                                          mul_add[2][164]<=((mult_out_20[164] + mult_out_21[164] + mult_out_22[164])%3329) ;
                                                                          mul_add[2][165]<=((mult_out_20[165] + mult_out_21[165] + mult_out_22[165])%3329) ;
                                                                          mul_add[2][166]<=((mult_out_20[166] + mult_out_21[166] + mult_out_22[166])%3329) ;
                                                                          mul_add[2][167]<=((mult_out_20[167] + mult_out_21[167] + mult_out_22[167])%3329) ;
                                                                          mul_add[2][168]<=((mult_out_20[168] + mult_out_21[168] + mult_out_22[168])%3329) ;
                                                                          mul_add[2][169]<=((mult_out_20[169] + mult_out_21[169] + mult_out_22[169])%3329) ;
                                                                          mul_add[2][170]<=((mult_out_20[170] + mult_out_21[170] + mult_out_22[170])%3329) ;
                                                                          mul_add[2][171]<=((mult_out_20[171] + mult_out_21[171] + mult_out_22[171])%3329) ;
                                                                          mul_add[2][172]<=((mult_out_20[172] + mult_out_21[172] + mult_out_22[172])%3329) ;
                                                                          mul_add[2][173]<=((mult_out_20[173] + mult_out_21[173] + mult_out_22[173])%3329) ;
                                                                          mul_add[2][174]<=((mult_out_20[174] + mult_out_21[174] + mult_out_22[174])%3329) ;
                                                                          mul_add[2][175]<=((mult_out_20[175] + mult_out_21[175] + mult_out_22[175])%3329) ;
                                                                          mul_add[2][176]<=((mult_out_20[176] + mult_out_21[176] + mult_out_22[176])%3329) ;
                                                                          mul_add[2][177]<=((mult_out_20[177] + mult_out_21[177] + mult_out_22[177])%3329) ;
                                                                          mul_add[2][178]<=((mult_out_20[178] + mult_out_21[178] + mult_out_22[178])%3329) ;
                                                                          mul_add[2][179]<=((mult_out_20[179] + mult_out_21[179] + mult_out_22[179])%3329) ;
                                                                          mul_add[2][180]<=((mult_out_20[180] + mult_out_21[180] + mult_out_22[180])%3329) ;
                                                                          mul_add[2][181]<=((mult_out_20[181] + mult_out_21[181] + mult_out_22[181])%3329) ;
                                                                          mul_add[2][182]<=((mult_out_20[182] + mult_out_21[182] + mult_out_22[182])%3329) ;
                                                                          mul_add[2][183]<=((mult_out_20[183] + mult_out_21[183] + mult_out_22[183])%3329) ;
                                                                          mul_add[2][184]<=((mult_out_20[184] + mult_out_21[184] + mult_out_22[184])%3329) ;
                                                                          mul_add[2][185]<=((mult_out_20[185] + mult_out_21[185] + mult_out_22[185])%3329) ;
                                                                          mul_add[2][186]<=((mult_out_20[186] + mult_out_21[186] + mult_out_22[186])%3329) ;
                                                                          mul_add[2][187]<=((mult_out_20[187] + mult_out_21[187] + mult_out_22[187])%3329) ;
                                                                          mul_add[2][188]<=((mult_out_20[188] + mult_out_21[188] + mult_out_22[188])%3329) ;
                                                                          mul_add[2][189]<=((mult_out_20[189] + mult_out_21[189] + mult_out_22[189])%3329) ;
                                                                          mul_add[2][190]<=((mult_out_20[190] + mult_out_21[190] + mult_out_22[190])%3329) ;
                                                                          mul_add[2][191]<=((mult_out_20[191] + mult_out_21[191] + mult_out_22[191])%3329) ;
                                                                          mul_add[2][192]<=((mult_out_20[192] + mult_out_21[192] + mult_out_22[192])%3329) ;
                                                                          mul_add[2][193]<=((mult_out_20[193] + mult_out_21[193] + mult_out_22[193])%3329) ;
                                                                          mul_add[2][194]<=((mult_out_20[194] + mult_out_21[194] + mult_out_22[194])%3329) ;
                                                                          mul_add[2][195]<=((mult_out_20[195] + mult_out_21[195] + mult_out_22[195])%3329) ;
                                                                          mul_add[2][196]<=((mult_out_20[196] + mult_out_21[196] + mult_out_22[196])%3329) ;
                                                                          mul_add[2][197]<=((mult_out_20[197] + mult_out_21[197] + mult_out_22[197])%3329) ;
                                                                          mul_add[2][198]<=((mult_out_20[198] + mult_out_21[198] + mult_out_22[198])%3329) ;
                                                                          mul_add[2][199]<=((mult_out_20[199] + mult_out_21[199] + mult_out_22[199])%3329) ;
                                                                          mul_add[2][200]<=((mult_out_20[200] + mult_out_21[200] + mult_out_22[200])%3329) ;
                                                                          mul_add[2][201]<=((mult_out_20[201] + mult_out_21[201] + mult_out_22[201])%3329) ;
                                                                          mul_add[2][202]<=((mult_out_20[202] + mult_out_21[202] + mult_out_22[202])%3329) ;
                                                                          mul_add[2][203]<=((mult_out_20[203] + mult_out_21[203] + mult_out_22[203])%3329) ;
                                                                          mul_add[2][204]<=((mult_out_20[204] + mult_out_21[204] + mult_out_22[204])%3329) ;
                                                                          mul_add[2][205]<=((mult_out_20[205] + mult_out_21[205] + mult_out_22[205])%3329) ;
                                                                          mul_add[2][206]<=((mult_out_20[206] + mult_out_21[206] + mult_out_22[206])%3329) ;
                                                                          mul_add[2][207]<=((mult_out_20[207] + mult_out_21[207] + mult_out_22[207])%3329) ;
                                                                          mul_add[2][208]<=((mult_out_20[208] + mult_out_21[208] + mult_out_22[208])%3329) ;
                                                                          mul_add[2][209]<=((mult_out_20[209] + mult_out_21[209] + mult_out_22[209])%3329) ;
                                                                          mul_add[2][210]<=((mult_out_20[210] + mult_out_21[210] + mult_out_22[210])%3329) ;
                                                                          mul_add[2][211]<=((mult_out_20[211] + mult_out_21[211] + mult_out_22[211])%3329) ;
                                                                          mul_add[2][212]<=((mult_out_20[212] + mult_out_21[212] + mult_out_22[212])%3329) ;
                                                                          mul_add[2][213]<=((mult_out_20[213] + mult_out_21[213] + mult_out_22[213])%3329) ;
                                                                          mul_add[2][214]<=((mult_out_20[214] + mult_out_21[214] + mult_out_22[214])%3329) ;
                                                                          mul_add[2][215]<=((mult_out_20[215] + mult_out_21[215] + mult_out_22[215])%3329) ;
                                                                          mul_add[2][216]<=((mult_out_20[216] + mult_out_21[216] + mult_out_22[216])%3329) ;
                                                                          mul_add[2][217]<=((mult_out_20[217] + mult_out_21[217] + mult_out_22[217])%3329) ;
                                                                          mul_add[2][218]<=((mult_out_20[218] + mult_out_21[218] + mult_out_22[218])%3329) ;
                                                                          mul_add[2][219]<=((mult_out_20[219] + mult_out_21[219] + mult_out_22[219])%3329) ;
                                                                          mul_add[2][220]<=((mult_out_20[220] + mult_out_21[220] + mult_out_22[220])%3329) ;
                                                                          mul_add[2][221]<=((mult_out_20[221] + mult_out_21[221] + mult_out_22[221])%3329) ;
                                                                          mul_add[2][222]<=((mult_out_20[222] + mult_out_21[222] + mult_out_22[222])%3329) ;
                                                                          mul_add[2][223]<=((mult_out_20[223] + mult_out_21[223] + mult_out_22[223])%3329) ;
                                                                          mul_add[2][224]<=((mult_out_20[224] + mult_out_21[224] + mult_out_22[224])%3329) ;
                                                                          mul_add[2][225]<=((mult_out_20[225] + mult_out_21[225] + mult_out_22[225])%3329) ;
                                                                          mul_add[2][226]<=((mult_out_20[226] + mult_out_21[226] + mult_out_22[226])%3329) ;
                                                                          mul_add[2][227]<=((mult_out_20[227] + mult_out_21[227] + mult_out_22[227])%3329) ;
                                                                          mul_add[2][228]<=((mult_out_20[228] + mult_out_21[228] + mult_out_22[228])%3329) ;
                                                                          mul_add[2][229]<=((mult_out_20[229] + mult_out_21[229] + mult_out_22[229])%3329) ;
                                                                          mul_add[2][230]<=((mult_out_20[230] + mult_out_21[230] + mult_out_22[230])%3329) ;
                                                                          mul_add[2][231]<=((mult_out_20[231] + mult_out_21[231] + mult_out_22[231])%3329) ;
                                                                          mul_add[2][232]<=((mult_out_20[232] + mult_out_21[232] + mult_out_22[232])%3329) ;
                                                                          mul_add[2][233]<=((mult_out_20[233] + mult_out_21[233] + mult_out_22[233])%3329) ;
                                                                          mul_add[2][234]<=((mult_out_20[234] + mult_out_21[234] + mult_out_22[234])%3329) ;
                                                                          mul_add[2][235]<=((mult_out_20[235] + mult_out_21[235] + mult_out_22[235])%3329) ;
                                                                          mul_add[2][236]<=((mult_out_20[236] + mult_out_21[236] + mult_out_22[236])%3329) ;
                                                                          mul_add[2][237]<=((mult_out_20[237] + mult_out_21[237] + mult_out_22[237])%3329) ;
                                                                          mul_add[2][238]<=((mult_out_20[238] + mult_out_21[238] + mult_out_22[238])%3329) ;
                                                                          mul_add[2][239]<=((mult_out_20[239] + mult_out_21[239] + mult_out_22[239])%3329) ;
                                                                          mul_add[2][240]<=((mult_out_20[240] + mult_out_21[240] + mult_out_22[240])%3329) ;
                                                                          mul_add[2][241]<=((mult_out_20[241] + mult_out_21[241] + mult_out_22[241])%3329) ;
                                                                          mul_add[2][242]<=((mult_out_20[242] + mult_out_21[242] + mult_out_22[242])%3329) ;
                                                                          mul_add[2][243]<=((mult_out_20[243] + mult_out_21[243] + mult_out_22[243])%3329) ;
                                                                          mul_add[2][244]<=((mult_out_20[244] + mult_out_21[244] + mult_out_22[244])%3329) ;
                                                                          mul_add[2][245]<=((mult_out_20[245] + mult_out_21[245] + mult_out_22[245])%3329) ;
                                                                          mul_add[2][246]<=((mult_out_20[246] + mult_out_21[246] + mult_out_22[246])%3329) ;
                                                                          mul_add[2][247]<=((mult_out_20[247] + mult_out_21[247] + mult_out_22[247])%3329) ;
                                                                          mul_add[2][248]<=((mult_out_20[248] + mult_out_21[248] + mult_out_22[248])%3329) ;
                                                                          mul_add[2][249]<=((mult_out_20[249] + mult_out_21[249] + mult_out_22[249])%3329) ;
                                                                          mul_add[2][250]<=((mult_out_20[250] + mult_out_21[250] + mult_out_22[250])%3329) ;
                                                                          mul_add[2][251]<=((mult_out_20[251] + mult_out_21[251] + mult_out_22[251])%3329) ;
                                                                          mul_add[2][252]<=((mult_out_20[252] + mult_out_21[252] + mult_out_22[252])%3329) ;
                                                                          mul_add[2][253]<=((mult_out_20[253] + mult_out_21[253] + mult_out_22[253])%3329) ;
                                                                          mul_add[2][254]<=((mult_out_20[254] + mult_out_21[254] + mult_out_22[254])%3329) ;
                                                                          mul_add[2][255]<=((mult_out_20[255] + mult_out_21[255] + mult_out_22[255])%3329) ;
                                                                
                                                                                          
                      multiply_ntts
                          mult_1 (
                              .clk(clk),
                              .reset(rst),
                              .f(T_hat_0),  // T_hat_0_16 is a 16-bit array
                              .g(y_ntt[0]),  // y_ntt_0_16 is now a 1D array
                              .zetas(zetas),
                              .h(mult_out_1),
                              .start(start_mul),
                              .done(done9_mul)
                          );
                      
                      multiply_ntts
                          mult_2 (
                              .clk(clk),
                              .reset(rst),
                              .f(T_hat_1),  // T_hat_1_16 is a 16-bit array
                              .g(y_ntt[1]),  // y_ntt_1_16 is now a 1D array
                              .zetas(zetas),
                              .h(mult_out_2),
                              .start(start_mul),
                              .done(done10_mul)
                          );
                      
                      multiply_ntts
                          mult_3 (
                              .clk(clk),
                              .reset(rst),
                              .f(T_hat_2),  
                              .g(y_ntt[2]),  
                              .zetas(zetas),
                              .h(mult_out_3),
                              .start(start_mul),
                              .done(done11_mul)
                          );
                          
//assign start_inverse = (done10_ntt && done11_ntt && done12_ntt );

////AT x Y inverse
////logic  [31:0] in_1 [256-1:0];

//inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_1 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_00),
//    .start_ntt(start_inverse),
//    .done_ntt(done10_ntt),
//    .f_hat(in_1)
//);

//inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_2 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_01),
//    .start_ntt(start_inverse),
//    .done_ntt(done11_ntt),
//    .f_hat(in_2)
//);

//inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_3 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_02),
//    .start_ntt(start_inverse),
//    .done_ntt(done12_ntt),
//    .f_hat(in_3)
//);


//inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_4 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_10),
//    .start_ntt(start_inverse),
//    .done_ntt(done4_ntt),
//    .f_hat(in_4)
//);

//inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_5 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_11),
//    .start_ntt(start_inverse),
//    .done_ntt(done5_ntt),
//    .f_hat(in_5)
//);

//inverse_ntt #(.N(NUM_COEFFS), .Q(3329), .F(3303)) inverse_6 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_12),
//    .start_ntt(start_inverse),
//    .done_ntt(done6_ntt),
//    .f_hat(in_6)
//);

//inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_7 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_20),
//    .start_ntt(start_inverse),
//    .done_ntt(done7_ntt),
//    .f_hat(in_7)
//);

//inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_8 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_21),
//    .start_ntt(start_inverse),
//    .done_ntt(done8_ntt),
//    .f_hat(in_8)
//);

//inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_9 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_22),
//    .start_ntt(start_inverse),
//    .done_ntt(done9_ntt),
//    .f_hat(in_9)
//);
  
//T hat x Y   
//logic  [31:0] v_in_1 [256-1:0];

//inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_v_1 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_1),
//    .start_ntt(start_inverse),
//    .done_ntt(done13_ntt),
//    .f_hat(v_in_1)
//);

//inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_v_2 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_2),
//    .start_ntt(start_inverse),
//    .done_ntt(done14_ntt),
//    .f_hat(v_in_2)
//);

//inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_v_3 (
//    .clk(clk),
//    .rst(rst),
//    .f(mult_out_3),
//    .start_ntt(start_inverse),
//    .done_ntt(done15_ntt),
//    .f_hat(v_in_3)
//);
 
//        logic [31:0] e1_ext [0:2][255:0];

//        assign e1_ext[0][0] = {30'd0, e1[0][0]};
//        assign e1_ext[0][1] = {30'd0, e1[0][1]};
//        assign e1_ext[0][2] = {30'd0, e1[0][2]};
//        assign e1_ext[0][3] = {30'd0, e1[0][3]};
//        assign e1_ext[0][4] = {30'd0, e1[0][4]};
//        assign e1_ext[0][5] = {30'd0, e1[0][5]};
//        assign e1_ext[0][6] = {30'd0, e1[0][6]};
//        assign e1_ext[0][7] = {30'd0, e1[0][7]};
//        assign e1_ext[0][8] = {30'd0, e1[0][8]};
//        assign e1_ext[0][9] = {30'd0, e1[0][9]};
//        assign e1_ext[0][10] = {30'd0, e1[0][10]};
//        assign e1_ext[0][11] = {30'd0, e1[0][11]};
//        assign e1_ext[0][12] = {30'd0, e1[0][12]};
//        assign e1_ext[0][13] = {30'd0, e1[0][13]};
//        assign e1_ext[0][14] = {30'd0, e1[0][14]};
//        assign e1_ext[0][15] = {30'd0, e1[0][15]};
//        assign e1_ext[0][16] = {30'd0, e1[0][16]};
//        assign e1_ext[0][17] = {30'd0, e1[0][17]};
//        assign e1_ext[0][18] = {30'd0, e1[0][18]};
//        assign e1_ext[0][19] = {30'd0, e1[0][19]};
//        assign e1_ext[0][20] = {30'd0, e1[0][20]};
//        assign e1_ext[0][21] = {30'd0, e1[0][21]};
//        assign e1_ext[0][22] = {30'd0, e1[0][22]};
//        assign e1_ext[0][23] = {30'd0, e1[0][23]};
//        assign e1_ext[0][24] = {30'd0, e1[0][24]};
//        assign e1_ext[0][25] = {30'd0, e1[0][25]};
//        assign e1_ext[0][26] = {30'd0, e1[0][26]};
//        assign e1_ext[0][27] = {30'd0, e1[0][27]};
//        assign e1_ext[0][28] = {30'd0, e1[0][28]};
//        assign e1_ext[0][29] = {30'd0, e1[0][29]};
//        assign e1_ext[0][30] = {30'd0, e1[0][30]};
//        assign e1_ext[0][31] = {30'd0, e1[0][31]};
//        assign e1_ext[0][32] = {30'd0, e1[0][32]};
//        assign e1_ext[0][33] = {30'd0, e1[0][33]};
//        assign e1_ext[0][34] = {30'd0, e1[0][34]};
//        assign e1_ext[0][35] = {30'd0, e1[0][35]};
//        assign e1_ext[0][36] = {30'd0, e1[0][36]};
//        assign e1_ext[0][37] = {30'd0, e1[0][37]};
//        assign e1_ext[0][38] = {30'd0, e1[0][38]};
//        assign e1_ext[0][39] = {30'd0, e1[0][39]};
//        assign e1_ext[0][40] = {30'd0, e1[0][40]};
//        assign e1_ext[0][41] = {30'd0, e1[0][41]};
//        assign e1_ext[0][42] = {30'd0, e1[0][42]};
//        assign e1_ext[0][43] = {30'd0, e1[0][43]};
//        assign e1_ext[0][44] = {30'd0, e1[0][44]};
//        assign e1_ext[0][45] = {30'd0, e1[0][45]};
//        assign e1_ext[0][46] = {30'd0, e1[0][46]};
//        assign e1_ext[0][47] = {30'd0, e1[0][47]};
//        assign e1_ext[0][48] = {30'd0, e1[0][48]};
//        assign e1_ext[0][49] = {30'd0, e1[0][49]};
//        assign e1_ext[0][50] = {30'd0, e1[0][50]};
//        assign e1_ext[0][51] = {30'd0, e1[0][51]};
//        assign e1_ext[0][52] = {30'd0, e1[0][52]};
//        assign e1_ext[0][53] = {30'd0, e1[0][53]};
//        assign e1_ext[0][54] = {30'd0, e1[0][54]};
//        assign e1_ext[0][55] = {30'd0, e1[0][55]};
//        assign e1_ext[0][56] = {30'd0, e1[0][56]};
//        assign e1_ext[0][57] = {30'd0, e1[0][57]};
//        assign e1_ext[0][58] = {30'd0, e1[0][58]};
//        assign e1_ext[0][59] = {30'd0, e1[0][59]};
//        assign e1_ext[0][60] = {30'd0, e1[0][60]};
//        assign e1_ext[0][61] = {30'd0, e1[0][61]};
//        assign e1_ext[0][62] = {30'd0, e1[0][62]};
//        assign e1_ext[0][63] = {30'd0, e1[0][63]};
//        assign e1_ext[0][64] = {30'd0, e1[0][64]};
//        assign e1_ext[0][65] = {30'd0, e1[0][65]};
//        assign e1_ext[0][66] = {30'd0, e1[0][66]};
//        assign e1_ext[0][67] = {30'd0, e1[0][67]};
//        assign e1_ext[0][68] = {30'd0, e1[0][68]};
//        assign e1_ext[0][69] = {30'd0, e1[0][69]};
//        assign e1_ext[0][70] = {30'd0, e1[0][70]};
//        assign e1_ext[0][71] = {30'd0, e1[0][71]};
//        assign e1_ext[0][72] = {30'd0, e1[0][72]};
//        assign e1_ext[0][73] = {30'd0, e1[0][73]};
//        assign e1_ext[0][74] = {30'd0, e1[0][74]};
//        assign e1_ext[0][75] = {30'd0, e1[0][75]};
//        assign e1_ext[0][76] = {30'd0, e1[0][76]};
//        assign e1_ext[0][77] = {30'd0, e1[0][77]};
//        assign e1_ext[0][78] = {30'd0, e1[0][78]};
//        assign e1_ext[0][79] = {30'd0, e1[0][79]};
//        assign e1_ext[0][80] = {30'd0, e1[0][80]};
//        assign e1_ext[0][81] = {30'd0, e1[0][81]};
//        assign e1_ext[0][82] = {30'd0, e1[0][82]};
//        assign e1_ext[0][83] = {30'd0, e1[0][83]};
//        assign e1_ext[0][84] = {30'd0, e1[0][84]};
//        assign e1_ext[0][85] = {30'd0, e1[0][85]};
//        assign e1_ext[0][86] = {30'd0, e1[0][86]};
//        assign e1_ext[0][87] = {30'd0, e1[0][87]};
//        assign e1_ext[0][88] = {30'd0, e1[0][88]};
//        assign e1_ext[0][89] = {30'd0, e1[0][89]};
//        assign e1_ext[0][90] = {30'd0, e1[0][90]};
//        assign e1_ext[0][91] = {30'd0, e1[0][91]};
//        assign e1_ext[0][92] = {30'd0, e1[0][92]};
//        assign e1_ext[0][93] = {30'd0, e1[0][93]};
//        assign e1_ext[0][94] = {30'd0, e1[0][94]};
//        assign e1_ext[0][95] = {30'd0, e1[0][95]};
//        assign e1_ext[0][96] = {30'd0, e1[0][96]};
//        assign e1_ext[0][97] = {30'd0, e1[0][97]};
//        assign e1_ext[0][98] = {30'd0, e1[0][98]};
//        assign e1_ext[0][99] = {30'd0, e1[0][99]};
//        assign e1_ext[0][100] = {30'd0, e1[0][100]};
//        assign e1_ext[0][101] = {30'd0, e1[0][101]};
//        assign e1_ext[0][102] = {30'd0, e1[0][102]};
//        assign e1_ext[0][103] = {30'd0, e1[0][103]};
//        assign e1_ext[0][104] = {30'd0, e1[0][104]};
//        assign e1_ext[0][105] = {30'd0, e1[0][105]};
//        assign e1_ext[0][106] = {30'd0, e1[0][106]};
//        assign e1_ext[0][107] = {30'd0, e1[0][107]};
//        assign e1_ext[0][108] = {30'd0, e1[0][108]};
//        assign e1_ext[0][109] = {30'd0, e1[0][109]};
//        assign e1_ext[0][110] = {30'd0, e1[0][110]};
//        assign e1_ext[0][111] = {30'd0, e1[0][111]};
//        assign e1_ext[0][112] = {30'd0, e1[0][112]};
//        assign e1_ext[0][113] = {30'd0, e1[0][113]};
//        assign e1_ext[0][114] = {30'd0, e1[0][114]};
//        assign e1_ext[0][115] = {30'd0, e1[0][115]};
//        assign e1_ext[0][116] = {30'd0, e1[0][116]};
//        assign e1_ext[0][117] = {30'd0, e1[0][117]};
//        assign e1_ext[0][118] = {30'd0, e1[0][118]};
//        assign e1_ext[0][119] = {30'd0, e1[0][119]};
//        assign e1_ext[0][120] = {30'd0, e1[0][120]};
//        assign e1_ext[0][121] = {30'd0, e1[0][121]};
//        assign e1_ext[0][122] = {30'd0, e1[0][122]};
//        assign e1_ext[0][123] = {30'd0, e1[0][123]};
//        assign e1_ext[0][124] = {30'd0, e1[0][124]};
//        assign e1_ext[0][125] = {30'd0, e1[0][125]};
//        assign e1_ext[0][126] = {30'd0, e1[0][126]};
//        assign e1_ext[0][127] = {30'd0, e1[0][127]};
//        assign e1_ext[0][128] = {30'd0, e1[0][128]};
//        assign e1_ext[0][129] = {30'd0, e1[0][129]};
//        assign e1_ext[0][130] = {30'd0, e1[0][130]};
//        assign e1_ext[0][131] = {30'd0, e1[0][131]};
//        assign e1_ext[0][132] = {30'd0, e1[0][132]};
//        assign e1_ext[0][133] = {30'd0, e1[0][133]};
//        assign e1_ext[0][134] = {30'd0, e1[0][134]};
//        assign e1_ext[0][135] = {30'd0, e1[0][135]};
//        assign e1_ext[0][136] = {30'd0, e1[0][136]};
//        assign e1_ext[0][137] = {30'd0, e1[0][137]};
//        assign e1_ext[0][138] = {30'd0, e1[0][138]};
//        assign e1_ext[0][139] = {30'd0, e1[0][139]};
//        assign e1_ext[0][140] = {30'd0, e1[0][140]};
//        assign e1_ext[0][141] = {30'd0, e1[0][141]};
//        assign e1_ext[0][142] = {30'd0, e1[0][142]};
//        assign e1_ext[0][143] = {30'd0, e1[0][143]};
//        assign e1_ext[0][144] = {30'd0, e1[0][144]};
//        assign e1_ext[0][145] = {30'd0, e1[0][145]};
//        assign e1_ext[0][146] = {30'd0, e1[0][146]};
//        assign e1_ext[0][147] = {30'd0, e1[0][147]};
//        assign e1_ext[0][148] = {30'd0, e1[0][148]};
//        assign e1_ext[0][149] = {30'd0, e1[0][149]};
//        assign e1_ext[0][150] = {30'd0, e1[0][150]};
//        assign e1_ext[0][151] = {30'd0, e1[0][151]};
//        assign e1_ext[0][152] = {30'd0, e1[0][152]};
//        assign e1_ext[0][153] = {30'd0, e1[0][153]};
//        assign e1_ext[0][154] = {30'd0, e1[0][154]};
//        assign e1_ext[0][155] = {30'd0, e1[0][155]};
//        assign e1_ext[0][156] = {30'd0, e1[0][156]};
//        assign e1_ext[0][157] = {30'd0, e1[0][157]};
//        assign e1_ext[0][158] = {30'd0, e1[0][158]};
//        assign e1_ext[0][159] = {30'd0, e1[0][159]};
//        assign e1_ext[0][160] = {30'd0, e1[0][160]};
//        assign e1_ext[0][161] = {30'd0, e1[0][161]};
//        assign e1_ext[0][162] = {30'd0, e1[0][162]};
//        assign e1_ext[0][163] = {30'd0, e1[0][163]};
//        assign e1_ext[0][164] = {30'd0, e1[0][164]};
//        assign e1_ext[0][165] = {30'd0, e1[0][165]};
//        assign e1_ext[0][166] = {30'd0, e1[0][166]};
//        assign e1_ext[0][167] = {30'd0, e1[0][167]};
//        assign e1_ext[0][168] = {30'd0, e1[0][168]};
//        assign e1_ext[0][169] = {30'd0, e1[0][169]};
//        assign e1_ext[0][170] = {30'd0, e1[0][170]};
//        assign e1_ext[0][171] = {30'd0, e1[0][171]};
//        assign e1_ext[0][172] = {30'd0, e1[0][172]};
//        assign e1_ext[0][173] = {30'd0, e1[0][173]};
//        assign e1_ext[0][174] = {30'd0, e1[0][174]};
//        assign e1_ext[0][175] = {30'd0, e1[0][175]};
//        assign e1_ext[0][176] = {30'd0, e1[0][176]};
//        assign e1_ext[0][177] = {30'd0, e1[0][177]};
//        assign e1_ext[0][178] = {30'd0, e1[0][178]};
//        assign e1_ext[0][179] = {30'd0, e1[0][179]};
//        assign e1_ext[0][180] = {30'd0, e1[0][180]};
//        assign e1_ext[0][181] = {30'd0, e1[0][181]};
//        assign e1_ext[0][182] = {30'd0, e1[0][182]};
//        assign e1_ext[0][183] = {30'd0, e1[0][183]};
//        assign e1_ext[0][184] = {30'd0, e1[0][184]};
//        assign e1_ext[0][185] = {30'd0, e1[0][185]};
//        assign e1_ext[0][186] = {30'd0, e1[0][186]};
//        assign e1_ext[0][187] = {30'd0, e1[0][187]};
//        assign e1_ext[0][188] = {30'd0, e1[0][188]};
//        assign e1_ext[0][189] = {30'd0, e1[0][189]};
//        assign e1_ext[0][190] = {30'd0, e1[0][190]};
//        assign e1_ext[0][191] = {30'd0, e1[0][191]};
//        assign e1_ext[0][192] = {30'd0, e1[0][192]};
//        assign e1_ext[0][193] = {30'd0, e1[0][193]};
//        assign e1_ext[0][194] = {30'd0, e1[0][194]};
//        assign e1_ext[0][195] = {30'd0, e1[0][195]};
//        assign e1_ext[0][196] = {30'd0, e1[0][196]};
//        assign e1_ext[0][197] = {30'd0, e1[0][197]};
//        assign e1_ext[0][198] = {30'd0, e1[0][198]};
//        assign e1_ext[0][199] = {30'd0, e1[0][199]};
//        assign e1_ext[0][200] = {30'd0, e1[0][200]};
//        assign e1_ext[0][201] = {30'd0, e1[0][201]};
//        assign e1_ext[0][202] = {30'd0, e1[0][202]};
//        assign e1_ext[0][203] = {30'd0, e1[0][203]};
//        assign e1_ext[0][204] = {30'd0, e1[0][204]};
//        assign e1_ext[0][205] = {30'd0, e1[0][205]};
//        assign e1_ext[0][206] = {30'd0, e1[0][206]};
//        assign e1_ext[0][207] = {30'd0, e1[0][207]};
//        assign e1_ext[0][208] = {30'd0, e1[0][208]};
//        assign e1_ext[0][209] = {30'd0, e1[0][209]};
//        assign e1_ext[0][210] = {30'd0, e1[0][210]};
//        assign e1_ext[0][211] = {30'd0, e1[0][211]};
//        assign e1_ext[0][212] = {30'd0, e1[0][212]};
//        assign e1_ext[0][213] = {30'd0, e1[0][213]};
//        assign e1_ext[0][214] = {30'd0, e1[0][214]};
//        assign e1_ext[0][215] = {30'd0, e1[0][215]};
//        assign e1_ext[0][216] = {30'd0, e1[0][216]};
//        assign e1_ext[0][217] = {30'd0, e1[0][217]};
//        assign e1_ext[0][218] = {30'd0, e1[0][218]};
//        assign e1_ext[0][219] = {30'd0, e1[0][219]};
//        assign e1_ext[0][220] = {30'd0, e1[0][220]};
//        assign e1_ext[0][221] = {30'd0, e1[0][221]};
//        assign e1_ext[0][222] = {30'd0, e1[0][222]};
//        assign e1_ext[0][223] = {30'd0, e1[0][223]};
//        assign e1_ext[0][224] = {30'd0, e1[0][224]};
//        assign e1_ext[0][225] = {30'd0, e1[0][225]};
//        assign e1_ext[0][226] = {30'd0, e1[0][226]};
//        assign e1_ext[0][227] = {30'd0, e1[0][227]};
//        assign e1_ext[0][228] = {30'd0, e1[0][228]};
//        assign e1_ext[0][229] = {30'd0, e1[0][229]};
//        assign e1_ext[0][230] = {30'd0, e1[0][230]};
//        assign e1_ext[0][231] = {30'd0, e1[0][231]};
//        assign e1_ext[0][232] = {30'd0, e1[0][232]};
//        assign e1_ext[0][233] = {30'd0, e1[0][233]};
//        assign e1_ext[0][234] = {30'd0, e1[0][234]};
//        assign e1_ext[0][235] = {30'd0, e1[0][235]};
//        assign e1_ext[0][236] = {30'd0, e1[0][236]};
//        assign e1_ext[0][237] = {30'd0, e1[0][237]};
//        assign e1_ext[0][238] = {30'd0, e1[0][238]};
//        assign e1_ext[0][239] = {30'd0, e1[0][239]};
//        assign e1_ext[0][240] = {30'd0, e1[0][240]};
//        assign e1_ext[0][241] = {30'd0, e1[0][241]};
//        assign e1_ext[0][242] = {30'd0, e1[0][242]};
//        assign e1_ext[0][243] = {30'd0, e1[0][243]};
//        assign e1_ext[0][244] = {30'd0, e1[0][244]};
//        assign e1_ext[0][245] = {30'd0, e1[0][245]};
//        assign e1_ext[0][246] = {30'd0, e1[0][246]};
//        assign e1_ext[0][247] = {30'd0, e1[0][247]};
//        assign e1_ext[0][248] = {30'd0, e1[0][248]};
//        assign e1_ext[0][249] = {30'd0, e1[0][249]};
//        assign e1_ext[0][250] = {30'd0, e1[0][250]};
//        assign e1_ext[0][251] = {30'd0, e1[0][251]};
//        assign e1_ext[0][252] = {30'd0, e1[0][252]};
//        assign e1_ext[0][253] = {30'd0, e1[0][253]};
//        assign e1_ext[0][254] = {30'd0, e1[0][254]};
//        assign e1_ext[0][255] = {30'd0, e1[0][255]};
//        assign e1_ext[1][0] = {30'd0, e1[1][0]};
//        assign e1_ext[1][1] = {30'd0, e1[1][1]};
//        assign e1_ext[1][2] = {30'd0, e1[1][2]};
//        assign e1_ext[1][3] = {30'd0, e1[1][3]};
////        assign e1_ext[1][4] = {30'd0, e1[1][4]};
//        assign e1_ext[1][5] = {30'd0, e1[1][5]};
//        assign e1_ext[1][6] = {30'd0, e1[1][6]};
//        assign e1_ext[1][7] = {30'd0, e1[1][7]};
//        assign e1_ext[1][8] = {30'd0, e1[1][8]};
//        assign e1_ext[1][9] = {30'd0, e1[1][9]};
//        assign e1_ext[1][10] = {30'd0, e1[1][10]};
//        assign e1_ext[1][11] = {30'd0, e1[1][11]};
//        assign e1_ext[1][12] = {30'd0, e1[1][12]};
//        assign e1_ext[1][13] = {30'd0, e1[1][13]};
//        assign e1_ext[1][14] = {30'd0, e1[1][14]};
//        assign e1_ext[1][15] = {30'd0, e1[1][15]};
//        assign e1_ext[1][16] = {30'd0, e1[1][16]};
//        assign e1_ext[1][17] = {30'd0, e1[1][17]};
//        assign e1_ext[1][18] = {30'd0, e1[1][18]};
//        assign e1_ext[1][19] = {30'd0, e1[1][19]};
//        assign e1_ext[1][20] = {30'd0, e1[1][20]};
//        assign e1_ext[1][21] = {30'd0, e1[1][21]};
//        assign e1_ext[1][22] = {30'd0, e1[1][22]};
//        assign e1_ext[1][23] = {30'd0, e1[1][23]};
//        assign e1_ext[1][24] = {30'd0, e1[1][24]};
//        assign e1_ext[1][25] = {30'd0, e1[1][25]};
//        assign e1_ext[1][26] = {30'd0, e1[1][26]};
//        assign e1_ext[1][27] = {30'd0, e1[1][27]};
//        assign e1_ext[1][28] = {30'd0, e1[1][28]};
//        assign e1_ext[1][29] = {30'd0, e1[1][29]};
//        assign e1_ext[1][30] = {30'd0, e1[1][30]};
//        assign e1_ext[1][31] = {30'd0, e1[1][31]};
//        assign e1_ext[1][32] = {30'd0, e1[1][32]};
//        assign e1_ext[1][33] = {30'd0, e1[1][33]};
//        assign e1_ext[1][34] = {30'd0, e1[1][34]};
//        assign e1_ext[1][35] = {30'd0, e1[1][35]};
//        assign e1_ext[1][36] = {30'd0, e1[1][36]};
//        assign e1_ext[1][37] = {30'd0, e1[1][37]};
//        assign e1_ext[1][38] = {30'd0, e1[1][38]};
//        assign e1_ext[1][39] = {30'd0, e1[1][39]};
//        assign e1_ext[1][40] = {30'd0, e1[1][40]};
//        assign e1_ext[1][41] = {30'd0, e1[1][41]};
//        assign e1_ext[1][42] = {30'd0, e1[1][42]};
//        assign e1_ext[1][43] = {30'd0, e1[1][43]};
//        assign e1_ext[1][44] = {30'd0, e1[1][44]};
//        assign e1_ext[1][45] = {30'd0, e1[1][45]};
//        assign e1_ext[1][46] = {30'd0, e1[1][46]};
//        assign e1_ext[1][47] = {30'd0, e1[1][47]};
//        assign e1_ext[1][48] = {30'd0, e1[1][48]};
//        assign e1_ext[1][49] = {30'd0, e1[1][49]};
//        assign e1_ext[1][50] = {30'd0, e1[1][50]};
//        assign e1_ext[1][51] = {30'd0, e1[1][51]};
//        assign e1_ext[1][52] = {30'd0, e1[1][52]};
//        assign e1_ext[1][53] = {30'd0, e1[1][53]};
//        assign e1_ext[1][54] = {30'd0, e1[1][54]};
//        assign e1_ext[1][55] = {30'd0, e1[1][55]};
//        assign e1_ext[1][56] = {30'd0, e1[1][56]};
//        assign e1_ext[1][57] = {30'd0, e1[1][57]};
//        assign e1_ext[1][58] = {30'd0, e1[1][58]};
//        assign e1_ext[1][59] = {30'd0, e1[1][59]};
//        assign e1_ext[1][60] = {30'd0, e1[1][60]};
//        assign e1_ext[1][61] = {30'd0, e1[1][61]};
//        assign e1_ext[1][62] = {30'd0, e1[1][62]};
//        assign e1_ext[1][63] = {30'd0, e1[1][63]};
//        assign e1_ext[1][64] = {30'd0, e1[1][64]};
//        assign e1_ext[1][65] = {30'd0, e1[1][65]};
//        assign e1_ext[1][66] = {30'd0, e1[1][66]};
//        assign e1_ext[1][67] = {30'd0, e1[1][67]};
//        assign e1_ext[1][68] = {30'd0, e1[1][68]};
//        assign e1_ext[1][69] = {30'd0, e1[1][69]};
//        assign e1_ext[1][70] = {30'd0, e1[1][70]};
//        assign e1_ext[1][71] = {30'd0, e1[1][71]};
//        assign e1_ext[1][72] = {30'd0, e1[1][72]};
//        assign e1_ext[1][73] = {30'd0, e1[1][73]};
//        assign e1_ext[1][74] = {30'd0, e1[1][74]};
//        assign e1_ext[1][75] = {30'd0, e1[1][75]};
//        assign e1_ext[1][76] = {30'd0, e1[1][76]};
//        assign e1_ext[1][77] = {30'd0, e1[1][77]};
//        assign e1_ext[1][78] = {30'd0, e1[1][78]};
//        assign e1_ext[1][79] = {30'd0, e1[1][79]};
//        assign e1_ext[1][80] = {30'd0, e1[1][80]};
//        assign e1_ext[1][81] = {30'd0, e1[1][81]};
//        assign e1_ext[1][82] = {30'd0, e1[1][82]};
//        assign e1_ext[1][83] = {30'd0, e1[1][83]};
//        assign e1_ext[1][84] = {30'd0, e1[1][84]};
//        assign e1_ext[1][85] = {30'd0, e1[1][85]};
//        assign e1_ext[1][86] = {30'd0, e1[1][86]};
//        assign e1_ext[1][87] = {30'd0, e1[1][87]};
//        assign e1_ext[1][88] = {30'd0, e1[1][88]};
//        assign e1_ext[1][89] = {30'd0, e1[1][89]};
//        assign e1_ext[1][90] = {30'd0, e1[1][90]};
//        assign e1_ext[1][91] = {30'd0, e1[1][91]};
//        assign e1_ext[1][92] = {30'd0, e1[1][92]};
//        assign e1_ext[1][93] = {30'd0, e1[1][93]};
//        assign e1_ext[1][94] = {30'd0, e1[1][94]};
//        assign e1_ext[1][95] = {30'd0, e1[1][95]};
//        assign e1_ext[1][96] = {30'd0, e1[1][96]};
//        assign e1_ext[1][97] = {30'd0, e1[1][97]};
//        assign e1_ext[1][98] = {30'd0, e1[1][98]};
//        assign e1_ext[1][99] = {30'd0, e1[1][99]};
//        assign e1_ext[1][100] = {30'd0, e1[1][100]};
//        assign e1_ext[1][101] = {30'd0, e1[1][101]};
//        assign e1_ext[1][102] = {30'd0, e1[1][102]};
//        assign e1_ext[1][103] = {30'd0, e1[1][103]};
//        assign e1_ext[1][104] = {30'd0, e1[1][104]};
//        assign e1_ext[1][105] = {30'd0, e1[1][105]};
//        assign e1_ext[1][106] = {30'd0, e1[1][106]};
//        assign e1_ext[1][107] = {30'd0, e1[1][107]};
//        assign e1_ext[1][108] = {30'd0, e1[1][108]};
//        assign e1_ext[1][109] = {30'd0, e1[1][109]};
//        assign e1_ext[1][110] = {30'd0, e1[1][110]};
//        assign e1_ext[1][111] = {30'd0, e1[1][111]};
//        assign e1_ext[1][112] = {30'd0, e1[1][112]};
//        assign e1_ext[1][113] = {30'd0, e1[1][113]};
//        assign e1_ext[1][114] = {30'd0, e1[1][114]};
//        assign e1_ext[1][115] = {30'd0, e1[1][115]};
//        assign e1_ext[1][116] = {30'd0, e1[1][116]};
//        assign e1_ext[1][117] = {30'd0, e1[1][117]};
//        assign e1_ext[1][118] = {30'd0, e1[1][118]};
//        assign e1_ext[1][119] = {30'd0, e1[1][119]};
//        assign e1_ext[1][120] = {30'd0, e1[1][120]};
//        assign e1_ext[1][121] = {30'd0, e1[1][121]};
//        assign e1_ext[1][122] = {30'd0, e1[1][122]};
//        assign e1_ext[1][123] = {30'd0, e1[1][123]};
//        assign e1_ext[1][124] = {30'd0, e1[1][124]};
//        assign e1_ext[1][125] = {30'd0, e1[1][125]};
//        assign e1_ext[1][126] = {30'd0, e1[1][126]};
//        assign e1_ext[1][127] = {30'd0, e1[1][127]};
//        assign e1_ext[1][128] = {30'd0, e1[1][128]};
//        assign e1_ext[1][129] = {30'd0, e1[1][129]};
//        assign e1_ext[1][130] = {30'd0, e1[1][130]};
//        assign e1_ext[1][131] = {30'd0, e1[1][131]};
//        assign e1_ext[1][132] = {30'd0, e1[1][132]};
//        assign e1_ext[1][133] = {30'd0, e1[1][133]};
//        assign e1_ext[1][134] = {30'd0, e1[1][134]};
//        assign e1_ext[1][135] = {30'd0, e1[1][135]};
//        assign e1_ext[1][136] = {30'd0, e1[1][136]};
//        assign e1_ext[1][137] = {30'd0, e1[1][137]};
//        assign e1_ext[1][138] = {30'd0, e1[1][138]};
//        assign e1_ext[1][139] = {30'd0, e1[1][139]};
//        assign e1_ext[1][140] = {30'd0, e1[1][140]};
//        assign e1_ext[1][141] = {30'd0, e1[1][141]};
//        assign e1_ext[1][142] = {30'd0, e1[1][142]};
//        assign e1_ext[1][143] = {30'd0, e1[1][143]};
//        assign e1_ext[1][144] = {30'd0, e1[1][144]};
//        assign e1_ext[1][145] = {30'd0, e1[1][145]};
//        assign e1_ext[1][146] = {30'd0, e1[1][146]};
//        assign e1_ext[1][147] = {30'd0, e1[1][147]};
//        assign e1_ext[1][148] = {30'd0, e1[1][148]};
//        assign e1_ext[1][149] = {30'd0, e1[1][149]};
//        assign e1_ext[1][150] = {30'd0, e1[1][150]};
//        assign e1_ext[1][151] = {30'd0, e1[1][151]};
//        assign e1_ext[1][152] = {30'd0, e1[1][152]};
//        assign e1_ext[1][153] = {30'd0, e1[1][153]};
//        assign e1_ext[1][154] = {30'd0, e1[1][154]};
//        assign e1_ext[1][155] = {30'd0, e1[1][155]};
//        assign e1_ext[1][156] = {30'd0, e1[1][156]};
//        assign e1_ext[1][157] = {30'd0, e1[1][157]};
//        assign e1_ext[1][158] = {30'd0, e1[1][158]};
//        assign e1_ext[1][159] = {30'd0, e1[1][159]};
//        assign e1_ext[1][160] = {30'd0, e1[1][160]};
//        assign e1_ext[1][161] = {30'd0, e1[1][161]};
//        assign e1_ext[1][162] = {30'd0, e1[1][162]};
//        assign e1_ext[1][163] = {30'd0, e1[1][163]};
//        assign e1_ext[1][164] = {30'd0, e1[1][164]};
//        assign e1_ext[1][165] = {30'd0, e1[1][165]};
//        assign e1_ext[1][166] = {30'd0, e1[1][166]};
//        assign e1_ext[1][167] = {30'd0, e1[1][167]};
//        assign e1_ext[1][168] = {30'd0, e1[1][168]};
//        assign e1_ext[1][169] = {30'd0, e1[1][169]};
//        assign e1_ext[1][170] = {30'd0, e1[1][170]};
//        assign e1_ext[1][171] = {30'd0, e1[1][171]};
//        assign e1_ext[1][172] = {30'd0, e1[1][172]};
//        assign e1_ext[1][173] = {30'd0, e1[1][173]};
//        assign e1_ext[1][174] = {30'd0, e1[1][174]};
//        assign e1_ext[1][175] = {30'd0, e1[1][175]};
//        assign e1_ext[1][176] = {30'd0, e1[1][176]};
//        assign e1_ext[1][177] = {30'd0, e1[1][177]};
//        assign e1_ext[1][178] = {30'd0, e1[1][178]};
//        assign e1_ext[1][179] = {30'd0, e1[1][179]};
//        assign e1_ext[1][180] = {30'd0, e1[1][180]};
//        assign e1_ext[1][181] = {30'd0, e1[1][181]};
//        assign e1_ext[1][182] = {30'd0, e1[1][182]};
//        assign e1_ext[1][183] = {30'd0, e1[1][183]};
//        assign e1_ext[1][184] = {30'd0, e1[1][184]};
//        assign e1_ext[1][185] = {30'd0, e1[1][185]};
//        assign e1_ext[1][186] = {30'd0, e1[1][186]};
//        assign e1_ext[1][187] = {30'd0, e1[1][187]};
//        assign e1_ext[1][188] = {30'd0, e1[1][188]};
//        assign e1_ext[1][189] = {30'd0, e1[1][189]};
//        assign e1_ext[1][190] = {30'd0, e1[1][190]};
//        assign e1_ext[1][191] = {30'd0, e1[1][191]};
//        assign e1_ext[1][192] = {30'd0, e1[1][192]};
//        assign e1_ext[1][193] = {30'd0, e1[1][193]};
//        assign e1_ext[1][194] = {30'd0, e1[1][194]};
//        assign e1_ext[1][195] = {30'd0, e1[1][195]};
//        assign e1_ext[1][196] = {30'd0, e1[1][196]};
//        assign e1_ext[1][197] = {30'd0, e1[1][197]};
//        assign e1_ext[1][198] = {30'd0, e1[1][198]};
//        assign e1_ext[1][199] = {30'd0, e1[1][199]};
//        assign e1_ext[1][200] = {30'd0, e1[1][200]};
//        assign e1_ext[1][201] = {30'd0, e1[1][201]};
//        assign e1_ext[1][202] = {30'd0, e1[1][202]};
//        assign e1_ext[1][203] = {30'd0, e1[1][203]};
//        assign e1_ext[1][204] = {30'd0, e1[1][204]};
//        assign e1_ext[1][205] = {30'd0, e1[1][205]};
//        assign e1_ext[1][206] = {30'd0, e1[1][206]};
//        assign e1_ext[1][207] = {30'd0, e1[1][207]};
//        assign e1_ext[1][208] = {30'd0, e1[1][208]};
//        assign e1_ext[1][209] = {30'd0, e1[1][209]};
//        assign e1_ext[1][210] = {30'd0, e1[1][210]};
//        assign e1_ext[1][211] = {30'd0, e1[1][211]};
//        assign e1_ext[1][212] = {30'd0, e1[1][212]};
//        assign e1_ext[1][213] = {30'd0, e1[1][213]};
//        assign e1_ext[1][214] = {30'd0, e1[1][214]};
//        assign e1_ext[1][215] = {30'd0, e1[1][215]};
//        assign e1_ext[1][216] = {30'd0, e1[1][216]};
//        assign e1_ext[1][217] = {30'd0, e1[1][217]};
//        assign e1_ext[1][218] = {30'd0, e1[1][218]};
//        assign e1_ext[1][219] = {30'd0, e1[1][219]};
//        assign e1_ext[1][220] = {30'd0, e1[1][220]};
//        assign e1_ext[1][221] = {30'd0, e1[1][221]};
//        assign e1_ext[1][222] = {30'd0, e1[1][222]};
//        assign e1_ext[1][223] = {30'd0, e1[1][223]};
//        assign e1_ext[1][224] = {30'd0, e1[1][224]};
//        assign e1_ext[1][225] = {30'd0, e1[1][225]};
//        assign e1_ext[1][226] = {30'd0, e1[1][226]};
//        assign e1_ext[1][227] = {30'd0, e1[1][227]};
//        assign e1_ext[1][228] = {30'd0, e1[1][228]};
//        assign e1_ext[1][229] = {30'd0, e1[1][229]};
//        assign e1_ext[1][230] = {30'd0, e1[1][230]};
//        assign e1_ext[1][231] = {30'd0, e1[1][231]};
//        assign e1_ext[1][232] = {30'd0, e1[1][232]};
//        assign e1_ext[1][233] = {30'd0, e1[1][233]};
//        assign e1_ext[1][234] = {30'd0, e1[1][234]};
//        assign e1_ext[1][235] = {30'd0, e1[1][235]};
//        assign e1_ext[1][236] = {30'd0, e1[1][236]};
//        assign e1_ext[1][237] = {30'd0, e1[1][237]};
//        assign e1_ext[1][238] = {30'd0, e1[1][238]};
//        assign e1_ext[1][239] = {30'd0, e1[1][239]};
//        assign e1_ext[1][240] = {30'd0, e1[1][240]};
//        assign e1_ext[1][241] = {30'd0, e1[1][241]};
//        assign e1_ext[1][242] = {30'd0, e1[1][242]};
//        assign e1_ext[1][243] = {30'd0, e1[1][243]};
//        assign e1_ext[1][244] = {30'd0, e1[1][244]};
//        assign e1_ext[1][245] = {30'd0, e1[1][245]};
//        assign e1_ext[1][246] = {30'd0, e1[1][246]};
//        assign e1_ext[1][247] = {30'd0, e1[1][247]};
//        assign e1_ext[1][248] = {30'd0, e1[1][248]};
//        assign e1_ext[1][249] = {30'd0, e1[1][249]};
//        assign e1_ext[1][250] = {30'd0, e1[1][250]};
//        assign e1_ext[1][251] = {30'd0, e1[1][251]};
//        assign e1_ext[1][252] = {30'd0, e1[1][252]};
//        assign e1_ext[1][253] = {30'd0, e1[1][253]};
//        assign e1_ext[1][254] = {30'd0, e1[1][254]};
//        assign e1_ext[1][255] = {30'd0, e1[1][255]};
//        assign e1_ext[2][0] = {30'd0, e1[2][0]};
//        assign e1_ext[2][1] = {30'd0, e1[2][1]};
//        assign e1_ext[2][2] = {30'd0, e1[2][2]};
//        assign e1_ext[2][3] = {30'd0, e1[2][3]};
//        assign e1_ext[2][4] = {30'd0, e1[2][4]};
//        assign e1_ext[2][5] = {30'd0, e1[2][5]};
//        assign e1_ext[2][6] = {30'd0, e1[2][6]};
//        assign e1_ext[2][7] = {30'd0, e1[2][7]};
//        assign e1_ext[2][8] = {30'd0, e1[2][8]};
//        assign e1_ext[2][9] = {30'd0, e1[2][9]};
//        assign e1_ext[2][10] = {30'd0, e1[2][10]};
//        assign e1_ext[2][11] = {30'd0, e1[2][11]};
//        assign e1_ext[2][12] = {30'd0, e1[2][12]};
//        assign e1_ext[2][13] = {30'd0, e1[2][13]};
//        assign e1_ext[2][14] = {30'd0, e1[2][14]};
//        assign e1_ext[2][15] = {30'd0, e1[2][15]};
//        assign e1_ext[2][16] = {30'd0, e1[2][16]};
//        assign e1_ext[2][17] = {30'd0, e1[2][17]};
//        assign e1_ext[2][18] = {30'd0, e1[2][18]};
//        assign e1_ext[2][19] = {30'd0, e1[2][19]};
//        assign e1_ext[2][20] = {30'd0, e1[2][20]};
//        assign e1_ext[2][21] = {30'd0, e1[2][21]};
//        assign e1_ext[2][22] = {30'd0, e1[2][22]};
//        assign e1_ext[2][23] = {30'd0, e1[2][23]};
//        assign e1_ext[2][24] = {30'd0, e1[2][24]};
//        assign e1_ext[2][25] = {30'd0, e1[2][25]};
//        assign e1_ext[2][26] = {30'd0, e1[2][26]};
//        assign e1_ext[2][27] = {30'd0, e1[2][27]};
//        assign e1_ext[2][28] = {30'd0, e1[2][28]};
//        assign e1_ext[2][29] = {30'd0, e1[2][29]};
//        assign e1_ext[2][30] = {30'd0, e1[2][30]};
//        assign e1_ext[2][31] = {30'd0, e1[2][31]};
//        assign e1_ext[2][32] = {30'd0, e1[2][32]};
//        assign e1_ext[2][33] = {30'd0, e1[2][33]};
//        assign e1_ext[2][34] = {30'd0, e1[2][34]};
//        assign e1_ext[2][35] = {30'd0, e1[2][35]};
//        assign e1_ext[2][36] = {30'd0, e1[2][36]};
//        assign e1_ext[2][37] = {30'd0, e1[2][37]};
//        assign e1_ext[2][38] = {30'd0, e1[2][38]};
//        assign e1_ext[2][39] = {30'd0, e1[2][39]};
//        assign e1_ext[2][40] = {30'd0, e1[2][40]};
//        assign e1_ext[2][41] = {30'd0, e1[2][41]};
//        assign e1_ext[2][42] = {30'd0, e1[2][42]};
//        assign e1_ext[2][43] = {30'd0, e1[2][43]};
//        assign e1_ext[2][44] = {30'd0, e1[2][44]};
//        assign e1_ext[2][45] = {30'd0, e1[2][45]};
//        assign e1_ext[2][46] = {30'd0, e1[2][46]};
//        assign e1_ext[2][47] = {30'd0, e1[2][47]};
//        assign e1_ext[2][48] = {30'd0, e1[2][48]};
//        assign e1_ext[2][49] = {30'd0, e1[2][49]};
//        assign e1_ext[2][50] = {30'd0, e1[2][50]};
//        assign e1_ext[2][51] = {30'd0, e1[2][51]};
//        assign e1_ext[2][52] = {30'd0, e1[2][52]};
//        assign e1_ext[2][53] = {30'd0, e1[2][53]};
//        assign e1_ext[2][54] = {30'd0, e1[2][54]};
//        assign e1_ext[2][55] = {30'd0, e1[2][55]};
//        assign e1_ext[2][56] = {30'd0, e1[2][56]};
//        assign e1_ext[2][57] = {30'd0, e1[2][57]};
//        assign e1_ext[2][58] = {30'd0, e1[2][58]};
//        assign e1_ext[2][59] = {30'd0, e1[2][59]};
//        assign e1_ext[2][60] = {30'd0, e1[2][60]};
//        assign e1_ext[2][61] = {30'd0, e1[2][61]};
//        assign e1_ext[2][62] = {30'd0, e1[2][62]};
//        assign e1_ext[2][63] = {30'd0, e1[2][63]};
//        assign e1_ext[2][64] = {30'd0, e1[2][64]};
//        assign e1_ext[2][65] = {30'd0, e1[2][65]};
//        assign e1_ext[2][66] = {30'd0, e1[2][66]};
//        assign e1_ext[2][67] = {30'd0, e1[2][67]};
//        assign e1_ext[2][68] = {30'd0, e1[2][68]};
//        assign e1_ext[2][69] = {30'd0, e1[2][69]};
//        assign e1_ext[2][70] = {30'd0, e1[2][70]};
//        assign e1_ext[2][71] = {30'd0, e1[2][71]};
//        assign e1_ext[2][72] = {30'd0, e1[2][72]};
//        assign e1_ext[2][73] = {30'd0, e1[2][73]};
//        assign e1_ext[2][74] = {30'd0, e1[2][74]};
//        assign e1_ext[2][75] = {30'd0, e1[2][75]};
//        assign e1_ext[2][76] = {30'd0, e1[2][76]};
//        assign e1_ext[2][77] = {30'd0, e1[2][77]};
//        assign e1_ext[2][78] = {30'd0, e1[2][78]};
//        assign e1_ext[2][79] = {30'd0, e1[2][79]};
//        assign e1_ext[2][80] = {30'd0, e1[2][80]};
//        assign e1_ext[2][81] = {30'd0, e1[2][81]};
//        assign e1_ext[2][82] = {30'd0, e1[2][82]};
//        assign e1_ext[2][83] = {30'd0, e1[2][83]};
//        assign e1_ext[2][84] = {30'd0, e1[2][84]};
//        assign e1_ext[2][85] = {30'd0, e1[2][85]};
//        assign e1_ext[2][86] = {30'd0, e1[2][86]};
//        assign e1_ext[2][87] = {30'd0, e1[2][87]};
//        assign e1_ext[2][88] = {30'd0, e1[2][88]};
//        assign e1_ext[2][89] = {30'd0, e1[2][89]};
//        assign e1_ext[2][90] = {30'd0, e1[2][90]};
//        assign e1_ext[2][91] = {30'd0, e1[2][91]};
//        assign e1_ext[2][92] = {30'd0, e1[2][92]};
//        assign e1_ext[2][93] = {30'd0, e1[2][93]};
//        assign e1_ext[2][94] = {30'd0, e1[2][94]};
//        assign e1_ext[2][95] = {30'd0, e1[2][95]};
//        assign e1_ext[2][96] = {30'd0, e1[2][96]};
//        assign e1_ext[2][97] = {30'd0, e1[2][97]};
//        assign e1_ext[2][98] = {30'd0, e1[2][98]};
//        assign e1_ext[2][99] = {30'd0, e1[2][99]};
//        assign e1_ext[2][100] = {30'd0, e1[2][100]};
//        assign e1_ext[2][101] = {30'd0, e1[2][101]};
//        assign e1_ext[2][102] = {30'd0, e1[2][102]};
//        assign e1_ext[2][103] = {30'd0, e1[2][103]};
//        assign e1_ext[2][104] = {30'd0, e1[2][104]};
//        assign e1_ext[2][105] = {30'd0, e1[2][105]};
//        assign e1_ext[2][106] = {30'd0, e1[2][106]};
//        assign e1_ext[2][107] = {30'd0, e1[2][107]};
//        assign e1_ext[2][108] = {30'd0, e1[2][108]};
//        assign e1_ext[2][109] = {30'd0, e1[2][109]};
//        assign e1_ext[2][110] = {30'd0, e1[2][110]};
//        assign e1_ext[2][111] = {30'd0, e1[2][111]};
//        assign e1_ext[2][112] = {30'd0, e1[2][112]};
//        assign e1_ext[2][113] = {30'd0, e1[2][113]};
//        assign e1_ext[2][114] = {30'd0, e1[2][114]};
//        assign e1_ext[2][115] = {30'd0, e1[2][115]};
//        assign e1_ext[2][116] = {30'd0, e1[2][116]};
//        assign e1_ext[2][117] = {30'd0, e1[2][117]};
//        assign e1_ext[2][118] = {30'd0, e1[2][118]};
//        assign e1_ext[2][119] = {30'd0, e1[2][119]};
//        assign e1_ext[2][120] = {30'd0, e1[2][120]};
//        assign e1_ext[2][121] = {30'd0, e1[2][121]};
//        assign e1_ext[2][122] = {30'd0, e1[2][122]};
//        assign e1_ext[2][123] = {30'd0, e1[2][123]};
//        assign e1_ext[2][124] = {30'd0, e1[2][124]};
//        assign e1_ext[2][125] = {30'd0, e1[2][125]};
//        assign e1_ext[2][126] = {30'd0, e1[2][126]};
//        assign e1_ext[2][127] = {30'd0, e1[2][127]};
//        assign e1_ext[2][128] = {30'd0, e1[2][128]};
//        assign e1_ext[2][129] = {30'd0, e1[2][129]};
//        assign e1_ext[2][130] = {30'd0, e1[2][130]};
//        assign e1_ext[2][131] = {30'd0, e1[2][131]};
//        assign e1_ext[2][132] = {30'd0, e1[2][132]};
//        assign e1_ext[2][133] = {30'd0, e1[2][133]};
//        assign e1_ext[2][134] = {30'd0, e1[2][134]};
//        assign e1_ext[2][135] = {30'd0, e1[2][135]};
//        assign e1_ext[2][136] = {30'd0, e1[2][136]};
//        assign e1_ext[2][137] = {30'd0, e1[2][137]};
//        assign e1_ext[2][138] = {30'd0, e1[2][138]};
//        assign e1_ext[2][139] = {30'd0, e1[2][139]};
//        assign e1_ext[2][140] = {30'd0, e1[2][140]};
//        assign e1_ext[2][141] = {30'd0, e1[2][141]};
//        assign e1_ext[2][142] = {30'd0, e1[2][142]};
//        assign e1_ext[2][143] = {30'd0, e1[2][143]};
//        assign e1_ext[2][144] = {30'd0, e1[2][144]};
//        assign e1_ext[2][145] = {30'd0, e1[2][145]};
//        assign e1_ext[2][146] = {30'd0, e1[2][146]};
//        assign e1_ext[2][147] = {30'd0, e1[2][147]};
//        assign e1_ext[2][148] = {30'd0, e1[2][148]};
//        assign e1_ext[2][149] = {30'd0, e1[2][149]};
//        assign e1_ext[2][150] = {30'd0, e1[2][150]};
//        assign e1_ext[2][151] = {30'd0, e1[2][151]};
//        assign e1_ext[2][152] = {30'd0, e1[2][152]};
//        assign e1_ext[2][153] = {30'd0, e1[2][153]};
//        assign e1_ext[2][154] = {30'd0, e1[2][154]};
//        assign e1_ext[2][155] = {30'd0, e1[2][155]};
//        assign e1_ext[2][156] = {30'd0, e1[2][156]};
//        assign e1_ext[2][157] = {30'd0, e1[2][157]};
//        assign e1_ext[2][158] = {30'd0, e1[2][158]};
//        assign e1_ext[2][159] = {30'd0, e1[2][159]};
//        assign e1_ext[2][160] = {30'd0, e1[2][160]};
//        assign e1_ext[2][161] = {30'd0, e1[2][161]};
//        assign e1_ext[2][162] = {30'd0, e1[2][162]};
//        assign e1_ext[2][163] = {30'd0, e1[2][163]};
//        assign e1_ext[2][164] = {30'd0, e1[2][164]};
//        assign e1_ext[2][165] = {30'd0, e1[2][165]};
//        assign e1_ext[2][166] = {30'd0, e1[2][166]};
//        assign e1_ext[2][167] = {30'd0, e1[2][167]};
//        assign e1_ext[2][168] = {30'd0, e1[2][168]};
//        assign e1_ext[2][169] = {30'd0, e1[2][169]};
//        assign e1_ext[2][170] = {30'd0, e1[2][170]};
//        assign e1_ext[2][171] = {30'd0, e1[2][171]};
//        assign e1_ext[2][172] = {30'd0, e1[2][172]};
//        assign e1_ext[2][173] = {30'd0, e1[2][173]};
//        assign e1_ext[2][174] = {30'd0, e1[2][174]};
//        assign e1_ext[2][175] = {30'd0, e1[2][175]};
//        assign e1_ext[2][176] = {30'd0, e1[2][176]};
//        assign e1_ext[2][177] = {30'd0, e1[2][177]};
//        assign e1_ext[2][178] = {30'd0, e1[2][178]};
//        assign e1_ext[2][179] = {30'd0, e1[2][179]};
//        assign e1_ext[2][180] = {30'd0, e1[2][180]};
//        assign e1_ext[2][181] = {30'd0, e1[2][181]};
//        assign e1_ext[2][182] = {30'd0, e1[2][182]};
//        assign e1_ext[2][183] = {30'd0, e1[2][183]};
//        assign e1_ext[2][184] = {30'd0, e1[2][184]};
//        assign e1_ext[2][185] = {30'd0, e1[2][185]};
//        assign e1_ext[2][186] = {30'd0, e1[2][186]};
//        assign e1_ext[2][187] = {30'd0, e1[2][187]};
//        assign e1_ext[2][188] = {30'd0, e1[2][188]};
//        assign e1_ext[2][189] = {30'd0, e1[2][189]};
//        assign e1_ext[2][190] = {30'd0, e1[2][190]};
//        assign e1_ext[2][191] = {30'd0, e1[2][191]};
//        assign e1_ext[2][192] = {30'd0, e1[2][192]};
//        assign e1_ext[2][193] = {30'd0, e1[2][193]};
//        assign e1_ext[2][194] = {30'd0, e1[2][194]};
//        assign e1_ext[2][195] = {30'd0, e1[2][195]};
//        assign e1_ext[2][196] = {30'd0, e1[2][196]};
//        assign e1_ext[2][197] = {30'd0, e1[2][197]};
//        assign e1_ext[2][198] = {30'd0, e1[2][198]};
//        assign e1_ext[2][199] = {30'd0, e1[2][199]};
//        assign e1_ext[2][200] = {30'd0, e1[2][200]};
//        assign e1_ext[2][201] = {30'd0, e1[2][201]};
//        assign e1_ext[2][202] = {30'd0, e1[2][202]};
//        assign e1_ext[2][203] = {30'd0, e1[2][203]};
//        assign e1_ext[2][204] = {30'd0, e1[2][204]};
//        assign e1_ext[2][205] = {30'd0, e1[2][205]};
//        assign e1_ext[2][206] = {30'd0, e1[2][206]};
//        assign e1_ext[2][207] = {30'd0, e1[2][207]};
//        assign e1_ext[2][208] = {30'd0, e1[2][208]};
//        assign e1_ext[2][209] = {30'd0, e1[2][209]};
//        assign e1_ext[2][210] = {30'd0, e1[2][210]};
//        assign e1_ext[2][211] = {30'd0, e1[2][211]};
//        assign e1_ext[2][212] = {30'd0, e1[2][212]};
//        assign e1_ext[2][213] = {30'd0, e1[2][213]};
//        assign e1_ext[2][214] = {30'd0, e1[2][214]};
//        assign e1_ext[2][215] = {30'd0, e1[2][215]};
//        assign e1_ext[2][216] = {30'd0, e1[2][216]};
//        assign e1_ext[2][217] = {30'd0, e1[2][217]};
//        assign e1_ext[2][218] = {30'd0, e1[2][218]};
//        assign e1_ext[2][219] = {30'd0, e1[2][219]};
//        assign e1_ext[2][220] = {30'd0, e1[2][220]};
//        assign e1_ext[2][221] = {30'd0, e1[2][221]};
//        assign e1_ext[2][222] = {30'd0, e1[2][222]};
//        assign e1_ext[2][223] = {30'd0, e1[2][223]};
//        assign e1_ext[2][224] = {30'd0, e1[2][224]};
//        assign e1_ext[2][225] = {30'd0, e1[2][225]};
//        assign e1_ext[2][226] = {30'd0, e1[2][226]};
//        assign e1_ext[2][227] = {30'd0, e1[2][227]};
//        assign e1_ext[2][228] = {30'd0, e1[2][228]};
//        assign e1_ext[2][229] = {30'd0, e1[2][229]};
//        assign e1_ext[2][230] = {30'd0, e1[2][230]};
//        assign e1_ext[2][231] = {30'd0, e1[2][231]};
//        assign e1_ext[2][232] = {30'd0, e1[2][232]};
//        assign e1_ext[2][233] = {30'd0, e1[2][233]};
//        assign e1_ext[2][234] = {30'd0, e1[2][234]};
//        assign e1_ext[2][235] = {30'd0, e1[2][235]};
//        assign e1_ext[2][236] = {30'd0, e1[2][236]};
//        assign e1_ext[2][237] = {30'd0, e1[2][237]};
//        assign e1_ext[2][238] = {30'd0, e1[2][238]};
//        assign e1_ext[2][239] = {30'd0, e1[2][239]};
//        assign e1_ext[2][240] = {30'd0, e1[2][240]};
//        assign e1_ext[2][241] = {30'd0, e1[2][241]};
//        assign e1_ext[2][242] = {30'd0, e1[2][242]};
//        assign e1_ext[2][243] = {30'd0, e1[2][243]};
//        assign e1_ext[2][244] = {30'd0, e1[2][244]};
//        assign e1_ext[2][245] = {30'd0, e1[2][245]};
//        assign e1_ext[2][246] = {30'd0, e1[2][246]};
//        assign e1_ext[2][247] = {30'd0, e1[2][247]};
//        assign e1_ext[2][248] = {30'd0, e1[2][248]};
//        assign e1_ext[2][249] = {30'd0, e1[2][249]};
//        assign e1_ext[2][250] = {30'd0, e1[2][250]};
//        assign e1_ext[2][251] = {30'd0, e1[2][251]};
//        assign e1_ext[2][252] = {30'd0, e1[2][252]};
//        assign e1_ext[2][253] = {30'd0, e1[2][253]};
//        assign e1_ext[2][254] = {30'd0, e1[2][254]};
//        assign e1_ext[2][255] = {30'd0, e1[2][255]};
        
////u = NTT_inverse(At x Y) + e1

//   assign u_1[0] = in_1[0] + e1_ext[0][0];
//   assign u_2[0] = in_2[0] + e1_ext[0][0];
//   assign u_3[0] = in_3[0] + e1_ext[0][0];
//   assign u_4[0] = in_4[0] + e1_ext[1][0];
//   assign u_5[0] = in_5[0] + e1_ext[1][0];
//   assign u_6[0] = in_6[0] + e1_ext[1][0];
//   assign u_7[0] = in_7[0] + e1_ext[2][0];
//   assign u_8[0] = in_8[0] + e1_ext[2][0];
//   assign u_9[0] = in_9[0] + e1_ext[2][0];
//   assign u_1[1] = in_1[1] + e1_ext[0][1];
//   assign u_2[1] = in_2[1] + e1_ext[0][1];
//   assign u_3[1] = in_3[1] + e1_ext[0][1];
//   assign u_4[1] = in_4[1] + e1_ext[1][1];
//   assign u_5[1] = in_5[1] + e1_ext[1][1];
//   assign u_6[1] = in_6[1] + e1_ext[1][1];
//   assign u_7[1] = in_7[1] + e1_ext[2][1];
//   assign u_8[1] = in_8[1] + e1_ext[2][1];
//   assign u_9[1] = in_9[1] + e1_ext[2][1];
//   assign u_1[2] = in_1[2] + e1_ext[0][2];
//   assign u_2[2] = in_2[2] + e1_ext[0][2];
//   assign u_3[2] = in_3[2] + e1_ext[0][2];
//   assign u_4[2] = in_4[2] + e1_ext[1][2];
//   assign u_5[2] = in_5[2] + e1_ext[1][2];
//   assign u_6[2] = in_6[2] + e1_ext[1][2];
//   assign u_7[2] = in_7[2] + e1_ext[2][2];
//   assign u_8[2] = in_8[2] + e1_ext[2][2];
//   assign u_9[2] = in_9[2] + e1_ext[2][2];
//   assign u_1[3] = in_1[3] + e1_ext[0][3];
//   assign u_2[3] = in_2[3] + e1_ext[0][3];
//   assign u_3[3] = in_3[3] + e1_ext[0][3];
//   assign u_4[3] = in_4[3] + e1_ext[1][3];
//   assign u_5[3] = in_5[3] + e1_ext[1][3];
//   assign u_6[3] = in_6[3] + e1_ext[1][3];
//   assign u_7[3] = in_7[3] + e1_ext[2][3];
//   assign u_8[3] = in_8[3] + e1_ext[2][3];
//   assign u_9[3] = in_9[3] + e1_ext[2][3];
//   assign u_1[4] = in_1[4] + e1_ext[0][4];
//   assign u_2[4] = in_2[4] + e1_ext[0][4];
//   assign u_3[4] = in_3[4] + e1_ext[0][4];
//   assign u_4[4] = in_4[4] + e1_ext[1][4];
//   assign u_5[4] = in_5[4] + e1_ext[1][4];
//   assign u_6[4] = in_6[4] + e1_ext[1][4];
//   assign u_7[4] = in_7[4] + e1_ext[2][4];
//   assign u_8[4] = in_8[4] + e1_ext[2][4];
//   assign u_9[4] = in_9[4] + e1_ext[2][4];
//   assign u_1[5] = in_1[5] + e1_ext[0][5];
//   assign u_2[5] = in_2[5] + e1_ext[0][5];
//   assign u_3[5] = in_3[5] + e1_ext[0][5];
//   assign u_4[5] = in_4[5] + e1_ext[1][5];
//   assign u_5[5] = in_5[5] + e1_ext[1][5];
//   assign u_6[5] = in_6[5] + e1_ext[1][5];
//   assign u_7[5] = in_7[5] + e1_ext[2][5];
//   assign u_8[5] = in_8[5] + e1_ext[2][5];
//   assign u_9[5] = in_9[5] + e1_ext[2][5];
//   assign u_1[6] = in_1[6] + e1_ext[0][6];
//   assign u_2[6] = in_2[6] + e1_ext[0][6];
//   assign u_3[6] = in_3[6] + e1_ext[0][6];
//   assign u_4[6] = in_4[6] + e1_ext[1][6];
//   assign u_5[6] = in_5[6] + e1_ext[1][6];
//   assign u_6[6] = in_6[6] + e1_ext[1][6];
//   assign u_7[6] = in_7[6] + e1_ext[2][6];
//   assign u_8[6] = in_8[6] + e1_ext[2][6];
//   assign u_9[6] = in_9[6] + e1_ext[2][6];
//   assign u_1[7] = in_1[7] + e1_ext[0][7];
//   assign u_2[7] = in_2[7] + e1_ext[0][7];
//   assign u_3[7] = in_3[7] + e1_ext[0][7];
//   assign u_4[7] = in_4[7] + e1_ext[1][7];
//   assign u_5[7] = in_5[7] + e1_ext[1][7];
//   assign u_6[7] = in_6[7] + e1_ext[1][7];
//   assign u_7[7] = in_7[7] + e1_ext[2][7];
//   assign u_8[7] = in_8[7] + e1_ext[2][7];
//   assign u_9[7] = in_9[7] + e1_ext[2][7];
//   assign u_1[8] = in_1[8] + e1_ext[0][8];
//   assign u_2[8] = in_2[8] + e1_ext[0][8];
//   assign u_3[8] = in_3[8] + e1_ext[0][8];
//   assign u_4[8] = in_4[8] + e1_ext[1][8];
//   assign u_5[8] = in_5[8] + e1_ext[1][8];
//   assign u_6[8] = in_6[8] + e1_ext[1][8];
//   assign u_7[8] = in_7[8] + e1_ext[2][8];
//   assign u_8[8] = in_8[8] + e1_ext[2][8];
//   assign u_9[8] = in_9[8] + e1_ext[2][8];
//   assign u_1[9] = in_1[9] + e1_ext[0][9];
//   assign u_2[9] = in_2[9] + e1_ext[0][9];
//   assign u_3[9] = in_3[9] + e1_ext[0][9];
//   assign u_4[9] = in_4[9] + e1_ext[1][9];
//   assign u_5[9] = in_5[9] + e1_ext[1][9];
//   assign u_6[9] = in_6[9] + e1_ext[1][9];
//   assign u_7[9] = in_7[9] + e1_ext[2][9];
//   assign u_8[9] = in_8[9] + e1_ext[2][9];
//   assign u_9[9] = in_9[9] + e1_ext[2][9];
//   assign u_1[10] = in_1[10] + e1_ext[0][10];
//   assign u_2[10] = in_2[10] + e1_ext[0][10];
//   assign u_3[10] = in_3[10] + e1_ext[0][10];
//   assign u_4[10] = in_4[10] + e1_ext[1][10];
//   assign u_5[10] = in_5[10] + e1_ext[1][10];
//   assign u_6[10] = in_6[10] + e1_ext[1][10];
//   assign u_7[10] = in_7[10] + e1_ext[2][10];
//   assign u_8[10] = in_8[10] + e1_ext[2][10];
//   assign u_9[10] = in_9[10] + e1_ext[2][10];
//   assign u_1[11] = in_1[11] + e1_ext[0][11];
//   assign u_2[11] = in_2[11] + e1_ext[0][11];
//   assign u_3[11] = in_3[11] + e1_ext[0][11];
//   assign u_4[11] = in_4[11] + e1_ext[1][11];
//   assign u_5[11] = in_5[11] + e1_ext[1][11];
//   assign u_6[11] = in_6[11] + e1_ext[1][11];
//   assign u_7[11] = in_7[11] + e1_ext[2][11];
//   assign u_8[11] = in_8[11] + e1_ext[2][11];
//   assign u_9[11] = in_9[11] + e1_ext[2][11];
//   assign u_1[12] = in_1[12] + e1_ext[0][12];
//   assign u_2[12] = in_2[12] + e1_ext[0][12];
//   assign u_3[12] = in_3[12] + e1_ext[0][12];
//   assign u_4[12] = in_4[12] + e1_ext[1][12];
//   assign u_5[12] = in_5[12] + e1_ext[1][12];
//   assign u_6[12] = in_6[12] + e1_ext[1][12];
//   assign u_7[12] = in_7[12] + e1_ext[2][12];
//   assign u_8[12] = in_8[12] + e1_ext[2][12];
//   assign u_9[12] = in_9[12] + e1_ext[2][12];
//   assign u_1[13] = in_1[13] + e1_ext[0][13];
//   assign u_2[13] = in_2[13] + e1_ext[0][13];
//   assign u_3[13] = in_3[13] + e1_ext[0][13];
//   assign u_4[13] = in_4[13] + e1_ext[1][13];
//   assign u_5[13] = in_5[13] + e1_ext[1][13];
//   assign u_6[13] = in_6[13] + e1_ext[1][13];
//   assign u_7[13] = in_7[13] + e1_ext[2][13];
//   assign u_8[13] = in_8[13] + e1_ext[2][13];
//   assign u_9[13] = in_9[13] + e1_ext[2][13];
//   assign u_1[14] = in_1[14] + e1_ext[0][14];
//   assign u_2[14] = in_2[14] + e1_ext[0][14];
//   assign u_3[14] = in_3[14] + e1_ext[0][14];
//   assign u_4[14] = in_4[14] + e1_ext[1][14];
//   assign u_5[14] = in_5[14] + e1_ext[1][14];
//   assign u_6[14] = in_6[14] + e1_ext[1][14];
//   assign u_7[14] = in_7[14] + e1_ext[2][14];
//   assign u_8[14] = in_8[14] + e1_ext[2][14];
//   assign u_9[14] = in_9[14] + e1_ext[2][14];
//   assign u_1[15] = in_1[15] + e1_ext[0][15];
//   assign u_2[15] = in_2[15] + e1_ext[0][15];
//   assign u_3[15] = in_3[15] + e1_ext[0][15];
//   assign u_4[15] = in_4[15] + e1_ext[1][15];
//   assign u_5[15] = in_5[15] + e1_ext[1][15];
//   assign u_6[15] = in_6[15] + e1_ext[1][15];
//   assign u_7[15] = in_7[15] + e1_ext[2][15];
//   assign u_8[15] = in_8[15] + e1_ext[2][15];
//   assign u_9[15] = in_9[15] + e1_ext[2][15];
//   assign u_1[16] = in_1[16] + e1_ext[0][16];
//   assign u_2[16] = in_2[16] + e1_ext[0][16];
//   assign u_3[16] = in_3[16] + e1_ext[0][16];
//   assign u_4[16] = in_4[16] + e1_ext[1][16];
//   assign u_5[16] = in_5[16] + e1_ext[1][16];
//   assign u_6[16] = in_6[16] + e1_ext[1][16];
//   assign u_7[16] = in_7[16] + e1_ext[2][16];
//   assign u_8[16] = in_8[16] + e1_ext[2][16];
//   assign u_9[16] = in_9[16] + e1_ext[2][16];
//   assign u_1[17] = in_1[17] + e1_ext[0][17];
//   assign u_2[17] = in_2[17] + e1_ext[0][17];
//   assign u_3[17] = in_3[17] + e1_ext[0][17];
//   assign u_4[17] = in_4[17] + e1_ext[1][17];
//   assign u_5[17] = in_5[17] + e1_ext[1][17];
//   assign u_6[17] = in_6[17] + e1_ext[1][17];
//   assign u_7[17] = in_7[17] + e1_ext[2][17];
//   assign u_8[17] = in_8[17] + e1_ext[2][17];
//   assign u_9[17] = in_9[17] + e1_ext[2][17];
//   assign u_1[18] = in_1[18] + e1_ext[0][18];
//   assign u_2[18] = in_2[18] + e1_ext[0][18];
//   assign u_3[18] = in_3[18] + e1_ext[0][18];
//   assign u_4[18] = in_4[18] + e1_ext[1][18];
//   assign u_5[18] = in_5[18] + e1_ext[1][18];
//   assign u_6[18] = in_6[18] + e1_ext[1][18];
//   assign u_7[18] = in_7[18] + e1_ext[2][18];
//   assign u_8[18] = in_8[18] + e1_ext[2][18];
//   assign u_9[18] = in_9[18] + e1_ext[2][18];
//   assign u_1[19] = in_1[19] + e1_ext[0][19];
//   assign u_2[19] = in_2[19] + e1_ext[0][19];
//   assign u_3[19] = in_3[19] + e1_ext[0][19];
//   assign u_4[19] = in_4[19] + e1_ext[1][19];
//   assign u_5[19] = in_5[19] + e1_ext[1][19];
//   assign u_6[19] = in_6[19] + e1_ext[1][19];
//   assign u_7[19] = in_7[19] + e1_ext[2][19];
//   assign u_8[19] = in_8[19] + e1_ext[2][19];
//   assign u_9[19] = in_9[19] + e1_ext[2][19];
//   assign u_1[20] = in_1[20] + e1_ext[0][20];
//   assign u_2[20] = in_2[20] + e1_ext[0][20];
//   assign u_3[20] = in_3[20] + e1_ext[0][20];
//   assign u_4[20] = in_4[20] + e1_ext[1][20];
//   assign u_5[20] = in_5[20] + e1_ext[1][20];
//   assign u_6[20] = in_6[20] + e1_ext[1][20];
//   assign u_7[20] = in_7[20] + e1_ext[2][20];
//   assign u_8[20] = in_8[20] + e1_ext[2][20];
//   assign u_9[20] = in_9[20] + e1_ext[2][20];
//   assign u_1[21] = in_1[21] + e1_ext[0][21];
//   assign u_2[21] = in_2[21] + e1_ext[0][21];
//   assign u_3[21] = in_3[21] + e1_ext[0][21];
//   assign u_4[21] = in_4[21] + e1_ext[1][21];
//   assign u_5[21] = in_5[21] + e1_ext[1][21];
//   assign u_6[21] = in_6[21] + e1_ext[1][21];
//   assign u_7[21] = in_7[21] + e1_ext[2][21];
//   assign u_8[21] = in_8[21] + e1_ext[2][21];
//   assign u_9[21] = in_9[21] + e1_ext[2][21];
//   assign u_1[22] = in_1[22] + e1_ext[0][22];
//   assign u_2[22] = in_2[22] + e1_ext[0][22];
//   assign u_3[22] = in_3[22] + e1_ext[0][22];
//   assign u_4[22] = in_4[22] + e1_ext[1][22];
//   assign u_5[22] = in_5[22] + e1_ext[1][22];
//   assign u_6[22] = in_6[22] + e1_ext[1][22];
//   assign u_7[22] = in_7[22] + e1_ext[2][22];
//   assign u_8[22] = in_8[22] + e1_ext[2][22];
//   assign u_9[22] = in_9[22] + e1_ext[2][22];
//   assign u_1[23] = in_1[23] + e1_ext[0][23];
//   assign u_2[23] = in_2[23] + e1_ext[0][23];
//   assign u_3[23] = in_3[23] + e1_ext[0][23];
//   assign u_4[23] = in_4[23] + e1_ext[1][23];
//   assign u_5[23] = in_5[23] + e1_ext[1][23];
//   assign u_6[23] = in_6[23] + e1_ext[1][23];
//   assign u_7[23] = in_7[23] + e1_ext[2][23];
//   assign u_8[23] = in_8[23] + e1_ext[2][23];
//   assign u_9[23] = in_9[23] + e1_ext[2][23];
//   assign u_1[24] = in_1[24] + e1_ext[0][24];
//   assign u_2[24] = in_2[24] + e1_ext[0][24];
//   assign u_3[24] = in_3[24] + e1_ext[0][24];
//   assign u_4[24] = in_4[24] + e1_ext[1][24];
//   assign u_5[24] = in_5[24] + e1_ext[1][24];
//   assign u_6[24] = in_6[24] + e1_ext[1][24];
//   assign u_7[24] = in_7[24] + e1_ext[2][24];
//   assign u_8[24] = in_8[24] + e1_ext[2][24];
//   assign u_9[24] = in_9[24] + e1_ext[2][24];
//   assign u_1[25] = in_1[25] + e1_ext[0][25];
//   assign u_2[25] = in_2[25] + e1_ext[0][25];
//   assign u_3[25] = in_3[25] + e1_ext[0][25];
//   assign u_4[25] = in_4[25] + e1_ext[1][25];
//   assign u_5[25] = in_5[25] + e1_ext[1][25];
//   assign u_6[25] = in_6[25] + e1_ext[1][25];
//   assign u_7[25] = in_7[25] + e1_ext[2][25];
//   assign u_8[25] = in_8[25] + e1_ext[2][25];
//   assign u_9[25] = in_9[25] + e1_ext[2][25];
//   assign u_1[26] = in_1[26] + e1_ext[0][26];
//   assign u_2[26] = in_2[26] + e1_ext[0][26];
//   assign u_3[26] = in_3[26] + e1_ext[0][26];
//   assign u_4[26] = in_4[26] + e1_ext[1][26];
//   assign u_5[26] = in_5[26] + e1_ext[1][26];
//   assign u_6[26] = in_6[26] + e1_ext[1][26];
//   assign u_7[26] = in_7[26] + e1_ext[2][26];
//   assign u_8[26] = in_8[26] + e1_ext[2][26];
//   assign u_9[26] = in_9[26] + e1_ext[2][26];
//   assign u_1[27] = in_1[27] + e1_ext[0][27];
//   assign u_2[27] = in_2[27] + e1_ext[0][27];
//   assign u_3[27] = in_3[27] + e1_ext[0][27];
//   assign u_4[27] = in_4[27] + e1_ext[1][27];
//   assign u_5[27] = in_5[27] + e1_ext[1][27];
//   assign u_6[27] = in_6[27] + e1_ext[1][27];
//   assign u_7[27] = in_7[27] + e1_ext[2][27];
//   assign u_8[27] = in_8[27] + e1_ext[2][27];
//   assign u_9[27] = in_9[27] + e1_ext[2][27];
//   assign u_1[28] = in_1[28] + e1_ext[0][28];
//   assign u_2[28] = in_2[28] + e1_ext[0][28];
//   assign u_3[28] = in_3[28] + e1_ext[0][28];
//   assign u_4[28] = in_4[28] + e1_ext[1][28];
//   assign u_5[28] = in_5[28] + e1_ext[1][28];
//   assign u_6[28] = in_6[28] + e1_ext[1][28];
//   assign u_7[28] = in_7[28] + e1_ext[2][28];
//   assign u_8[28] = in_8[28] + e1_ext[2][28];
//   assign u_9[28] = in_9[28] + e1_ext[2][28];
//   assign u_1[29] = in_1[29] + e1_ext[0][29];
//   assign u_2[29] = in_2[29] + e1_ext[0][29];
//   assign u_3[29] = in_3[29] + e1_ext[0][29];
//   assign u_4[29] = in_4[29] + e1_ext[1][29];
//   assign u_5[29] = in_5[29] + e1_ext[1][29];
//   assign u_6[29] = in_6[29] + e1_ext[1][29];
//   assign u_7[29] = in_7[29] + e1_ext[2][29];
//   assign u_8[29] = in_8[29] + e1_ext[2][29];
//   assign u_9[29] = in_9[29] + e1_ext[2][29];
//   assign u_1[30] = in_1[30] + e1_ext[0][30];
//   assign u_2[30] = in_2[30] + e1_ext[0][30];
//   assign u_3[30] = in_3[30] + e1_ext[0][30];
//   assign u_4[30] = in_4[30] + e1_ext[1][30];
//   assign u_5[30] = in_5[30] + e1_ext[1][30];
//   assign u_6[30] = in_6[30] + e1_ext[1][30];
//   assign u_7[30] = in_7[30] + e1_ext[2][30];
//   assign u_8[30] = in_8[30] + e1_ext[2][30];
//   assign u_9[30] = in_9[30] + e1_ext[2][30];
//   assign u_1[31] = in_1[31] + e1_ext[0][31];
//   assign u_2[31] = in_2[31] + e1_ext[0][31];
//   assign u_3[31] = in_3[31] + e1_ext[0][31];
//   assign u_4[31] = in_4[31] + e1_ext[1][31];
//   assign u_5[31] = in_5[31] + e1_ext[1][31];
//   assign u_6[31] = in_6[31] + e1_ext[1][31];
//   assign u_7[31] = in_7[31] + e1_ext[2][31];
//   assign u_8[31] = in_8[31] + e1_ext[2][31];
//   assign u_9[31] = in_9[31] + e1_ext[2][31];
//   assign u_1[32] = in_1[32] + e1_ext[0][32];
//   assign u_2[32] = in_2[32] + e1_ext[0][32];
//   assign u_3[32] = in_3[32] + e1_ext[0][32];
//   assign u_4[32] = in_4[32] + e1_ext[1][32];
//   assign u_5[32] = in_5[32] + e1_ext[1][32];
//   assign u_6[32] = in_6[32] + e1_ext[1][32];
//   assign u_7[32] = in_7[32] + e1_ext[2][32];
//   assign u_8[32] = in_8[32] + e1_ext[2][32];
//   assign u_9[32] = in_9[32] + e1_ext[2][32];
//   assign u_1[33] = in_1[33] + e1_ext[0][33];
//   assign u_2[33] = in_2[33] + e1_ext[0][33];
//   assign u_3[33] = in_3[33] + e1_ext[0][33];
//   assign u_4[33] = in_4[33] + e1_ext[1][33];
//   assign u_5[33] = in_5[33] + e1_ext[1][33];
//   assign u_6[33] = in_6[33] + e1_ext[1][33];
//   assign u_7[33] = in_7[33] + e1_ext[2][33];
//   assign u_8[33] = in_8[33] + e1_ext[2][33];
//   assign u_9[33] = in_9[33] + e1_ext[2][33];
//   assign u_1[34] = in_1[34] + e1_ext[0][34];
//   assign u_2[34] = in_2[34] + e1_ext[0][34];
//   assign u_3[34] = in_3[34] + e1_ext[0][34];
//   assign u_4[34] = in_4[34] + e1_ext[1][34];
//   assign u_5[34] = in_5[34] + e1_ext[1][34];
//   assign u_6[34] = in_6[34] + e1_ext[1][34];
//   assign u_7[34] = in_7[34] + e1_ext[2][34];
//   assign u_8[34] = in_8[34] + e1_ext[2][34];
//   assign u_9[34] = in_9[34] + e1_ext[2][34];
//   assign u_1[35] = in_1[35] + e1_ext[0][35];
//   assign u_2[35] = in_2[35] + e1_ext[0][35];
//   assign u_3[35] = in_3[35] + e1_ext[0][35];
//   assign u_4[35] = in_4[35] + e1_ext[1][35];
//   assign u_5[35] = in_5[35] + e1_ext[1][35];
//   assign u_6[35] = in_6[35] + e1_ext[1][35];
//   assign u_7[35] = in_7[35] + e1_ext[2][35];
//   assign u_8[35] = in_8[35] + e1_ext[2][35];
//   assign u_9[35] = in_9[35] + e1_ext[2][35];
//   assign u_1[36] = in_1[36] + e1_ext[0][36];
//   assign u_2[36] = in_2[36] + e1_ext[0][36];
//   assign u_3[36] = in_3[36] + e1_ext[0][36];
//   assign u_4[36] = in_4[36] + e1_ext[1][36];
//   assign u_5[36] = in_5[36] + e1_ext[1][36];
//   assign u_6[36] = in_6[36] + e1_ext[1][36];
//   assign u_7[36] = in_7[36] + e1_ext[2][36];
//   assign u_8[36] = in_8[36] + e1_ext[2][36];
//   assign u_9[36] = in_9[36] + e1_ext[2][36];
//   assign u_1[37] = in_1[37] + e1_ext[0][37];
//   assign u_2[37] = in_2[37] + e1_ext[0][37];
//   assign u_3[37] = in_3[37] + e1_ext[0][37];
//   assign u_4[37] = in_4[37] + e1_ext[1][37];
//   assign u_5[37] = in_5[37] + e1_ext[1][37];
//   assign u_6[37] = in_6[37] + e1_ext[1][37];
//   assign u_7[37] = in_7[37] + e1_ext[2][37];
//   assign u_8[37] = in_8[37] + e1_ext[2][37];
//   assign u_9[37] = in_9[37] + e1_ext[2][37];
//   assign u_1[38] = in_1[38] + e1_ext[0][38];
//   assign u_2[38] = in_2[38] + e1_ext[0][38];
//   assign u_3[38] = in_3[38] + e1_ext[0][38];
//   assign u_4[38] = in_4[38] + e1_ext[1][38];
//   assign u_5[38] = in_5[38] + e1_ext[1][38];
//   assign u_6[38] = in_6[38] + e1_ext[1][38];
//   assign u_7[38] = in_7[38] + e1_ext[2][38];
//   assign u_8[38] = in_8[38] + e1_ext[2][38];
//   assign u_9[38] = in_9[38] + e1_ext[2][38];
//   assign u_1[39] = in_1[39] + e1_ext[0][39];
//   assign u_2[39] = in_2[39] + e1_ext[0][39];
//   assign u_3[39] = in_3[39] + e1_ext[0][39];
//   assign u_4[39] = in_4[39] + e1_ext[1][39];
//   assign u_5[39] = in_5[39] + e1_ext[1][39];
//   assign u_6[39] = in_6[39] + e1_ext[1][39];
//   assign u_7[39] = in_7[39] + e1_ext[2][39];
//   assign u_8[39] = in_8[39] + e1_ext[2][39];
//   assign u_9[39] = in_9[39] + e1_ext[2][39];
//   assign u_1[40] = in_1[40] + e1_ext[0][40];
//   assign u_2[40] = in_2[40] + e1_ext[0][40];
//   assign u_3[40] = in_3[40] + e1_ext[0][40];
//   assign u_4[40] = in_4[40] + e1_ext[1][40];
//   assign u_5[40] = in_5[40] + e1_ext[1][40];
//   assign u_6[40] = in_6[40] + e1_ext[1][40];
//   assign u_7[40] = in_7[40] + e1_ext[2][40];
//   assign u_8[40] = in_8[40] + e1_ext[2][40];
//   assign u_9[40] = in_9[40] + e1_ext[2][40];
//   assign u_1[41] = in_1[41] + e1_ext[0][41];
//   assign u_2[41] = in_2[41] + e1_ext[0][41];
//   assign u_3[41] = in_3[41] + e1_ext[0][41];
//   assign u_4[41] = in_4[41] + e1_ext[1][41];
//   assign u_5[41] = in_5[41] + e1_ext[1][41];
//   assign u_6[41] = in_6[41] + e1_ext[1][41];
//   assign u_7[41] = in_7[41] + e1_ext[2][41];
//   assign u_8[41] = in_8[41] + e1_ext[2][41];
//   assign u_9[41] = in_9[41] + e1_ext[2][41];
//   assign u_1[42] = in_1[42] + e1_ext[0][42];
//   assign u_2[42] = in_2[42] + e1_ext[0][42];
//   assign u_3[42] = in_3[42] + e1_ext[0][42];
//   assign u_4[42] = in_4[42] + e1_ext[1][42];
//   assign u_5[42] = in_5[42] + e1_ext[1][42];
//   assign u_6[42] = in_6[42] + e1_ext[1][42];
//   assign u_7[42] = in_7[42] + e1_ext[2][42];
//   assign u_8[42] = in_8[42] + e1_ext[2][42];
//   assign u_9[42] = in_9[42] + e1_ext[2][42];
//   assign u_1[43] = in_1[43] + e1_ext[0][43];
//   assign u_2[43] = in_2[43] + e1_ext[0][43];
//   assign u_3[43] = in_3[43] + e1_ext[0][43];
//   assign u_4[43] = in_4[43] + e1_ext[1][43];
//   assign u_5[43] = in_5[43] + e1_ext[1][43];
//   assign u_6[43] = in_6[43] + e1_ext[1][43];
//   assign u_7[43] = in_7[43] + e1_ext[2][43];
//   assign u_8[43] = in_8[43] + e1_ext[2][43];
//   assign u_9[43] = in_9[43] + e1_ext[2][43];
//   assign u_1[44] = in_1[44] + e1_ext[0][44];
//   assign u_2[44] = in_2[44] + e1_ext[0][44];
//   assign u_3[44] = in_3[44] + e1_ext[0][44];
//   assign u_4[44] = in_4[44] + e1_ext[1][44];
//   assign u_5[44] = in_5[44] + e1_ext[1][44];
//   assign u_6[44] = in_6[44] + e1_ext[1][44];
//   assign u_7[44] = in_7[44] + e1_ext[2][44];
//   assign u_8[44] = in_8[44] + e1_ext[2][44];
//   assign u_9[44] = in_9[44] + e1_ext[2][44];
//   assign u_1[45] = in_1[45] + e1_ext[0][45];
//   assign u_2[45] = in_2[45] + e1_ext[0][45];
//   assign u_3[45] = in_3[45] + e1_ext[0][45];
//   assign u_4[45] = in_4[45] + e1_ext[1][45];
//   assign u_5[45] = in_5[45] + e1_ext[1][45];
//   assign u_6[45] = in_6[45] + e1_ext[1][45];
//   assign u_7[45] = in_7[45] + e1_ext[2][45];
//   assign u_8[45] = in_8[45] + e1_ext[2][45];
//   assign u_9[45] = in_9[45] + e1_ext[2][45];
//   assign u_1[46] = in_1[46] + e1_ext[0][46];
//   assign u_2[46] = in_2[46] + e1_ext[0][46];
//   assign u_3[46] = in_3[46] + e1_ext[0][46];
//   assign u_4[46] = in_4[46] + e1_ext[1][46];
//   assign u_5[46] = in_5[46] + e1_ext[1][46];
//   assign u_6[46] = in_6[46] + e1_ext[1][46];
//   assign u_7[46] = in_7[46] + e1_ext[2][46];
//   assign u_8[46] = in_8[46] + e1_ext[2][46];
//   assign u_9[46] = in_9[46] + e1_ext[2][46];
//   assign u_1[47] = in_1[47] + e1_ext[0][47];
//   assign u_2[47] = in_2[47] + e1_ext[0][47];
//   assign u_3[47] = in_3[47] + e1_ext[0][47];
//   assign u_4[47] = in_4[47] + e1_ext[1][47];
//   assign u_5[47] = in_5[47] + e1_ext[1][47];
//   assign u_6[47] = in_6[47] + e1_ext[1][47];
//   assign u_7[47] = in_7[47] + e1_ext[2][47];
//   assign u_8[47] = in_8[47] + e1_ext[2][47];
//   assign u_9[47] = in_9[47] + e1_ext[2][47];
//   assign u_1[48] = in_1[48] + e1_ext[0][48];
//   assign u_2[48] = in_2[48] + e1_ext[0][48];
//   assign u_3[48] = in_3[48] + e1_ext[0][48];
//   assign u_4[48] = in_4[48] + e1_ext[1][48];
//   assign u_5[48] = in_5[48] + e1_ext[1][48];
//   assign u_6[48] = in_6[48] + e1_ext[1][48];
//   assign u_7[48] = in_7[48] + e1_ext[2][48];
//   assign u_8[48] = in_8[48] + e1_ext[2][48];
//   assign u_9[48] = in_9[48] + e1_ext[2][48];
//   assign u_1[49] = in_1[49] + e1_ext[0][49];
//   assign u_2[49] = in_2[49] + e1_ext[0][49];
//   assign u_3[49] = in_3[49] + e1_ext[0][49];
//   assign u_4[49] = in_4[49] + e1_ext[1][49];
//   assign u_5[49] = in_5[49] + e1_ext[1][49];
//   assign u_6[49] = in_6[49] + e1_ext[1][49];
//   assign u_7[49] = in_7[49] + e1_ext[2][49];
//   assign u_8[49] = in_8[49] + e1_ext[2][49];
//   assign u_9[49] = in_9[49] + e1_ext[2][49];
//   assign u_1[50] = in_1[50] + e1_ext[0][50];
//   assign u_2[50] = in_2[50] + e1_ext[0][50];
//   assign u_3[50] = in_3[50] + e1_ext[0][50];
//   assign u_4[50] = in_4[50] + e1_ext[1][50];
//   assign u_5[50] = in_5[50] + e1_ext[1][50];
//   assign u_6[50] = in_6[50] + e1_ext[1][50];
//   assign u_7[50] = in_7[50] + e1_ext[2][50];
//   assign u_8[50] = in_8[50] + e1_ext[2][50];
//   assign u_9[50] = in_9[50] + e1_ext[2][50];
//   assign u_1[51] = in_1[51] + e1_ext[0][51];
//   assign u_2[51] = in_2[51] + e1_ext[0][51];
//   assign u_3[51] = in_3[51] + e1_ext[0][51];
//   assign u_4[51] = in_4[51] + e1_ext[1][51];
//   assign u_5[51] = in_5[51] + e1_ext[1][51];
//   assign u_6[51] = in_6[51] + e1_ext[1][51];
//   assign u_7[51] = in_7[51] + e1_ext[2][51];
//   assign u_8[51] = in_8[51] + e1_ext[2][51];
//   assign u_9[51] = in_9[51] + e1_ext[2][51];
//   assign u_1[52] = in_1[52] + e1_ext[0][52];
//   assign u_2[52] = in_2[52] + e1_ext[0][52];
//   assign u_3[52] = in_3[52] + e1_ext[0][52];
//   assign u_4[52] = in_4[52] + e1_ext[1][52];
//   assign u_5[52] = in_5[52] + e1_ext[1][52];
//   assign u_6[52] = in_6[52] + e1_ext[1][52];
//   assign u_7[52] = in_7[52] + e1_ext[2][52];
//   assign u_8[52] = in_8[52] + e1_ext[2][52];
//   assign u_9[52] = in_9[52] + e1_ext[2][52];
//   assign u_1[53] = in_1[53] + e1_ext[0][53];
//   assign u_2[53] = in_2[53] + e1_ext[0][53];
//   assign u_3[53] = in_3[53] + e1_ext[0][53];
//   assign u_4[53] = in_4[53] + e1_ext[1][53];
//   assign u_5[53] = in_5[53] + e1_ext[1][53];
//   assign u_6[53] = in_6[53] + e1_ext[1][53];
//   assign u_7[53] = in_7[53] + e1_ext[2][53];
//   assign u_8[53] = in_8[53] + e1_ext[2][53];
//   assign u_9[53] = in_9[53] + e1_ext[2][53];
//   assign u_1[54] = in_1[54] + e1_ext[0][54];
//   assign u_2[54] = in_2[54] + e1_ext[0][54];
//   assign u_3[54] = in_3[54] + e1_ext[0][54];
//   assign u_4[54] = in_4[54] + e1_ext[1][54];
//   assign u_5[54] = in_5[54] + e1_ext[1][54];
//   assign u_6[54] = in_6[54] + e1_ext[1][54];
//   assign u_7[54] = in_7[54] + e1_ext[2][54];
//   assign u_8[54] = in_8[54] + e1_ext[2][54];
//   assign u_9[54] = in_9[54] + e1_ext[2][54];
//   assign u_1[55] = in_1[55] + e1_ext[0][55];
//   assign u_2[55] = in_2[55] + e1_ext[0][55];
//   assign u_3[55] = in_3[55] + e1_ext[0][55];
//   assign u_4[55] = in_4[55] + e1_ext[1][55];
//   assign u_5[55] = in_5[55] + e1_ext[1][55];
//   assign u_6[55] = in_6[55] + e1_ext[1][55];
//   assign u_7[55] = in_7[55] + e1_ext[2][55];
//   assign u_8[55] = in_8[55] + e1_ext[2][55];
//   assign u_9[55] = in_9[55] + e1_ext[2][55];
//   assign u_1[56] = in_1[56] + e1_ext[0][56];
//   assign u_2[56] = in_2[56] + e1_ext[0][56];
//   assign u_3[56] = in_3[56] + e1_ext[0][56];
//   assign u_4[56] = in_4[56] + e1_ext[1][56];
//   assign u_5[56] = in_5[56] + e1_ext[1][56];
//   assign u_6[56] = in_6[56] + e1_ext[1][56];
//   assign u_7[56] = in_7[56] + e1_ext[2][56];
//   assign u_8[56] = in_8[56] + e1_ext[2][56];
//   assign u_9[56] = in_9[56] + e1_ext[2][56];
//   assign u_1[57] = in_1[57] + e1_ext[0][57];
//   assign u_2[57] = in_2[57] + e1_ext[0][57];
//   assign u_3[57] = in_3[57] + e1_ext[0][57];
//   assign u_4[57] = in_4[57] + e1_ext[1][57];
//   assign u_5[57] = in_5[57] + e1_ext[1][57];
//   assign u_6[57] = in_6[57] + e1_ext[1][57];
//   assign u_7[57] = in_7[57] + e1_ext[2][57];
//   assign u_8[57] = in_8[57] + e1_ext[2][57];
//   assign u_9[57] = in_9[57] + e1_ext[2][57];
//   assign u_1[58] = in_1[58] + e1_ext[0][58];
//   assign u_2[58] = in_2[58] + e1_ext[0][58];
//   assign u_3[58] = in_3[58] + e1_ext[0][58];
//   assign u_4[58] = in_4[58] + e1_ext[1][58];
//   assign u_5[58] = in_5[58] + e1_ext[1][58];
//   assign u_6[58] = in_6[58] + e1_ext[1][58];
//   assign u_7[58] = in_7[58] + e1_ext[2][58];
//   assign u_8[58] = in_8[58] + e1_ext[2][58];
//   assign u_9[58] = in_9[58] + e1_ext[2][58];
//   assign u_1[59] = in_1[59] + e1_ext[0][59];
//   assign u_2[59] = in_2[59] + e1_ext[0][59];
//   assign u_3[59] = in_3[59] + e1_ext[0][59];
//   assign u_4[59] = in_4[59] + e1_ext[1][59];
//   assign u_5[59] = in_5[59] + e1_ext[1][59];
//   assign u_6[59] = in_6[59] + e1_ext[1][59];
//   assign u_7[59] = in_7[59] + e1_ext[2][59];
//   assign u_8[59] = in_8[59] + e1_ext[2][59];
//   assign u_9[59] = in_9[59] + e1_ext[2][59];
//   assign u_1[60] = in_1[60] + e1_ext[0][60];
//   assign u_2[60] = in_2[60] + e1_ext[0][60];
//   assign u_3[60] = in_3[60] + e1_ext[0][60];
//   assign u_4[60] = in_4[60] + e1_ext[1][60];
//   assign u_5[60] = in_5[60] + e1_ext[1][60];
//   assign u_6[60] = in_6[60] + e1_ext[1][60];
//   assign u_7[60] = in_7[60] + e1_ext[2][60];
//   assign u_8[60] = in_8[60] + e1_ext[2][60];
//   assign u_9[60] = in_9[60] + e1_ext[2][60];
//   assign u_1[61] = in_1[61] + e1_ext[0][61];
//   assign u_2[61] = in_2[61] + e1_ext[0][61];
//   assign u_3[61] = in_3[61] + e1_ext[0][61];
//   assign u_4[61] = in_4[61] + e1_ext[1][61];
//   assign u_5[61] = in_5[61] + e1_ext[1][61];
//   assign u_6[61] = in_6[61] + e1_ext[1][61];
//   assign u_7[61] = in_7[61] + e1_ext[2][61];
//   assign u_8[61] = in_8[61] + e1_ext[2][61];
//   assign u_9[61] = in_9[61] + e1_ext[2][61];
//   assign u_1[62] = in_1[62] + e1_ext[0][62];
//   assign u_2[62] = in_2[62] + e1_ext[0][62];
//   assign u_3[62] = in_3[62] + e1_ext[0][62];
//   assign u_4[62] = in_4[62] + e1_ext[1][62];
//   assign u_5[62] = in_5[62] + e1_ext[1][62];
//   assign u_6[62] = in_6[62] + e1_ext[1][62];
//   assign u_7[62] = in_7[62] + e1_ext[2][62];
//   assign u_8[62] = in_8[62] + e1_ext[2][62];
//   assign u_9[62] = in_9[62] + e1_ext[2][62];
//   assign u_1[63] = in_1[63] + e1_ext[0][63];
//   assign u_2[63] = in_2[63] + e1_ext[0][63];
//   assign u_3[63] = in_3[63] + e1_ext[0][63];
//   assign u_4[63] = in_4[63] + e1_ext[1][63];
//   assign u_5[63] = in_5[63] + e1_ext[1][63];
//   assign u_6[63] = in_6[63] + e1_ext[1][63];
//   assign u_7[63] = in_7[63] + e1_ext[2][63];
//   assign u_8[63] = in_8[63] + e1_ext[2][63];
//   assign u_9[63] = in_9[63] + e1_ext[2][63];
//   assign u_1[64] = in_1[64] + e1_ext[0][64];
//   assign u_2[64] = in_2[64] + e1_ext[0][64];
//   assign u_3[64] = in_3[64] + e1_ext[0][64];
//   assign u_4[64] = in_4[64] + e1_ext[1][64];
//   assign u_5[64] = in_5[64] + e1_ext[1][64];
//   assign u_6[64] = in_6[64] + e1_ext[1][64];
//   assign u_7[64] = in_7[64] + e1_ext[2][64];
//   assign u_8[64] = in_8[64] + e1_ext[2][64];
//   assign u_9[64] = in_9[64] + e1_ext[2][64];
//   assign u_1[65] = in_1[65] + e1_ext[0][65];
//   assign u_2[65] = in_2[65] + e1_ext[0][65];
//   assign u_3[65] = in_3[65] + e1_ext[0][65];
//   assign u_4[65] = in_4[65] + e1_ext[1][65];
//   assign u_5[65] = in_5[65] + e1_ext[1][65];
//   assign u_6[65] = in_6[65] + e1_ext[1][65];
//   assign u_7[65] = in_7[65] + e1_ext[2][65];
//   assign u_8[65] = in_8[65] + e1_ext[2][65];
//   assign u_9[65] = in_9[65] + e1_ext[2][65];
//   assign u_1[66] = in_1[66] + e1_ext[0][66];
//   assign u_2[66] = in_2[66] + e1_ext[0][66];
//   assign u_3[66] = in_3[66] + e1_ext[0][66];
//   assign u_4[66] = in_4[66] + e1_ext[1][66];
//   assign u_5[66] = in_5[66] + e1_ext[1][66];
//   assign u_6[66] = in_6[66] + e1_ext[1][66];
//   assign u_7[66] = in_7[66] + e1_ext[2][66];
//   assign u_8[66] = in_8[66] + e1_ext[2][66];
//   assign u_9[66] = in_9[66] + e1_ext[2][66];
//   assign u_1[67] = in_1[67] + e1_ext[0][67];
//   assign u_2[67] = in_2[67] + e1_ext[0][67];
//   assign u_3[67] = in_3[67] + e1_ext[0][67];
//   assign u_4[67] = in_4[67] + e1_ext[1][67];
//   assign u_5[67] = in_5[67] + e1_ext[1][67];
//   assign u_6[67] = in_6[67] + e1_ext[1][67];
//   assign u_7[67] = in_7[67] + e1_ext[2][67];
//   assign u_8[67] = in_8[67] + e1_ext[2][67];
//   assign u_9[67] = in_9[67] + e1_ext[2][67];
//   assign u_1[68] = in_1[68] + e1_ext[0][68];
//   assign u_2[68] = in_2[68] + e1_ext[0][68];
//   assign u_3[68] = in_3[68] + e1_ext[0][68];
//   assign u_4[68] = in_4[68] + e1_ext[1][68];
//   assign u_5[68] = in_5[68] + e1_ext[1][68];
//   assign u_6[68] = in_6[68] + e1_ext[1][68];
//   assign u_7[68] = in_7[68] + e1_ext[2][68];
//   assign u_8[68] = in_8[68] + e1_ext[2][68];
//   assign u_9[68] = in_9[68] + e1_ext[2][68];
//   assign u_1[69] = in_1[69] + e1_ext[0][69];
//   assign u_2[69] = in_2[69] + e1_ext[0][69];
//   assign u_3[69] = in_3[69] + e1_ext[0][69];
//   assign u_4[69] = in_4[69] + e1_ext[1][69];
//   assign u_5[69] = in_5[69] + e1_ext[1][69];
//   assign u_6[69] = in_6[69] + e1_ext[1][69];
//   assign u_7[69] = in_7[69] + e1_ext[2][69];
//   assign u_8[69] = in_8[69] + e1_ext[2][69];
//   assign u_9[69] = in_9[69] + e1_ext[2][69];
//   assign u_1[70] = in_1[70] + e1_ext[0][70];
//   assign u_2[70] = in_2[70] + e1_ext[0][70];
//   assign u_3[70] = in_3[70] + e1_ext[0][70];
//   assign u_4[70] = in_4[70] + e1_ext[1][70];
//   assign u_5[70] = in_5[70] + e1_ext[1][70];
//   assign u_6[70] = in_6[70] + e1_ext[1][70];
//   assign u_7[70] = in_7[70] + e1_ext[2][70];
//   assign u_8[70] = in_8[70] + e1_ext[2][70];
//   assign u_9[70] = in_9[70] + e1_ext[2][70];
//   assign u_1[71] = in_1[71] + e1_ext[0][71];
//   assign u_2[71] = in_2[71] + e1_ext[0][71];
//   assign u_3[71] = in_3[71] + e1_ext[0][71];
//   assign u_4[71] = in_4[71] + e1_ext[1][71];
//   assign u_5[71] = in_5[71] + e1_ext[1][71];
//   assign u_6[71] = in_6[71] + e1_ext[1][71];
//   assign u_7[71] = in_7[71] + e1_ext[2][71];
//   assign u_8[71] = in_8[71] + e1_ext[2][71];
//   assign u_9[71] = in_9[71] + e1_ext[2][71];
//   assign u_1[72] = in_1[72] + e1_ext[0][72];
//   assign u_2[72] = in_2[72] + e1_ext[0][72];
//   assign u_3[72] = in_3[72] + e1_ext[0][72];
//   assign u_4[72] = in_4[72] + e1_ext[1][72];
//   assign u_5[72] = in_5[72] + e1_ext[1][72];
//   assign u_6[72] = in_6[72] + e1_ext[1][72];
//   assign u_7[72] = in_7[72] + e1_ext[2][72];
//   assign u_8[72] = in_8[72] + e1_ext[2][72];
//   assign u_9[72] = in_9[72] + e1_ext[2][72];
//   assign u_1[73] = in_1[73] + e1_ext[0][73];
//   assign u_2[73] = in_2[73] + e1_ext[0][73];
//   assign u_3[73] = in_3[73] + e1_ext[0][73];
//   assign u_4[73] = in_4[73] + e1_ext[1][73];
//   assign u_5[73] = in_5[73] + e1_ext[1][73];
//   assign u_6[73] = in_6[73] + e1_ext[1][73];
//   assign u_7[73] = in_7[73] + e1_ext[2][73];
//   assign u_8[73] = in_8[73] + e1_ext[2][73];
//   assign u_9[73] = in_9[73] + e1_ext[2][73];
//   assign u_1[74] = in_1[74] + e1_ext[0][74];
//   assign u_2[74] = in_2[74] + e1_ext[0][74];
//   assign u_3[74] = in_3[74] + e1_ext[0][74];
//   assign u_4[74] = in_4[74] + e1_ext[1][74];
//   assign u_5[74] = in_5[74] + e1_ext[1][74];
//   assign u_6[74] = in_6[74] + e1_ext[1][74];
//   assign u_7[74] = in_7[74] + e1_ext[2][74];
//   assign u_8[74] = in_8[74] + e1_ext[2][74];
//   assign u_9[74] = in_9[74] + e1_ext[2][74];
//   assign u_1[75] = in_1[75] + e1_ext[0][75];
//   assign u_2[75] = in_2[75] + e1_ext[0][75];
//   assign u_3[75] = in_3[75] + e1_ext[0][75];
//   assign u_4[75] = in_4[75] + e1_ext[1][75];
//   assign u_5[75] = in_5[75] + e1_ext[1][75];
//   assign u_6[75] = in_6[75] + e1_ext[1][75];
//   assign u_7[75] = in_7[75] + e1_ext[2][75];
//   assign u_8[75] = in_8[75] + e1_ext[2][75];
//   assign u_9[75] = in_9[75] + e1_ext[2][75];
//   assign u_1[76] = in_1[76] + e1_ext[0][76];
//   assign u_2[76] = in_2[76] + e1_ext[0][76];
//   assign u_3[76] = in_3[76] + e1_ext[0][76];
//   assign u_4[76] = in_4[76] + e1_ext[1][76];
//   assign u_5[76] = in_5[76] + e1_ext[1][76];
//   assign u_6[76] = in_6[76] + e1_ext[1][76];
//   assign u_7[76] = in_7[76] + e1_ext[2][76];
//   assign u_8[76] = in_8[76] + e1_ext[2][76];
//   assign u_9[76] = in_9[76] + e1_ext[2][76];
//   assign u_1[77] = in_1[77] + e1_ext[0][77];
//   assign u_2[77] = in_2[77] + e1_ext[0][77];
//   assign u_3[77] = in_3[77] + e1_ext[0][77];
//   assign u_4[77] = in_4[77] + e1_ext[1][77];
//   assign u_5[77] = in_5[77] + e1_ext[1][77];
//   assign u_6[77] = in_6[77] + e1_ext[1][77];
//   assign u_7[77] = in_7[77] + e1_ext[2][77];
//   assign u_8[77] = in_8[77] + e1_ext[2][77];
//   assign u_9[77] = in_9[77] + e1_ext[2][77];
//   assign u_1[78] = in_1[78] + e1_ext[0][78];
//   assign u_2[78] = in_2[78] + e1_ext[0][78];
//   assign u_3[78] = in_3[78] + e1_ext[0][78];
//   assign u_4[78] = in_4[78] + e1_ext[1][78];
//   assign u_5[78] = in_5[78] + e1_ext[1][78];
//   assign u_6[78] = in_6[78] + e1_ext[1][78];
//   assign u_7[78] = in_7[78] + e1_ext[2][78];
//   assign u_8[78] = in_8[78] + e1_ext[2][78];
//   assign u_9[78] = in_9[78] + e1_ext[2][78];
//   assign u_1[79] = in_1[79] + e1_ext[0][79];
//   assign u_2[79] = in_2[79] + e1_ext[0][79];
//   assign u_3[79] = in_3[79] + e1_ext[0][79];
//   assign u_4[79] = in_4[79] + e1_ext[1][79];
//   assign u_5[79] = in_5[79] + e1_ext[1][79];
//   assign u_6[79] = in_6[79] + e1_ext[1][79];
//   assign u_7[79] = in_7[79] + e1_ext[2][79];
//   assign u_8[79] = in_8[79] + e1_ext[2][79];
//   assign u_9[79] = in_9[79] + e1_ext[2][79];
//   assign u_1[80] = in_1[80] + e1_ext[0][80];
//   assign u_2[80] = in_2[80] + e1_ext[0][80];
//   assign u_3[80] = in_3[80] + e1_ext[0][80];
//   assign u_4[80] = in_4[80] + e1_ext[1][80];
//   assign u_5[80] = in_5[80] + e1_ext[1][80];
//   assign u_6[80] = in_6[80] + e1_ext[1][80];
//   assign u_7[80] = in_7[80] + e1_ext[2][80];
//   assign u_8[80] = in_8[80] + e1_ext[2][80];
//   assign u_9[80] = in_9[80] + e1_ext[2][80];
//   assign u_1[81] = in_1[81] + e1_ext[0][81];
//   assign u_2[81] = in_2[81] + e1_ext[0][81];
//   assign u_3[81] = in_3[81] + e1_ext[0][81];
//   assign u_4[81] = in_4[81] + e1_ext[1][81];
//   assign u_5[81] = in_5[81] + e1_ext[1][81];
//   assign u_6[81] = in_6[81] + e1_ext[1][81];
//   assign u_7[81] = in_7[81] + e1_ext[2][81];
//   assign u_8[81] = in_8[81] + e1_ext[2][81];
//   assign u_9[81] = in_9[81] + e1_ext[2][81];
//   assign u_1[82] = in_1[82] + e1_ext[0][82];
//   assign u_2[82] = in_2[82] + e1_ext[0][82];
//   assign u_3[82] = in_3[82] + e1_ext[0][82];
//   assign u_4[82] = in_4[82] + e1_ext[1][82];
//   assign u_5[82] = in_5[82] + e1_ext[1][82];
//   assign u_6[82] = in_6[82] + e1_ext[1][82];
//   assign u_7[82] = in_7[82] + e1_ext[2][82];
//   assign u_8[82] = in_8[82] + e1_ext[2][82];
//   assign u_9[82] = in_9[82] + e1_ext[2][82];
//   assign u_1[83] = in_1[83] + e1_ext[0][83];
//   assign u_2[83] = in_2[83] + e1_ext[0][83];
//   assign u_3[83] = in_3[83] + e1_ext[0][83];
//   assign u_4[83] = in_4[83] + e1_ext[1][83];
//   assign u_5[83] = in_5[83] + e1_ext[1][83];
//   assign u_6[83] = in_6[83] + e1_ext[1][83];
//   assign u_7[83] = in_7[83] + e1_ext[2][83];
//   assign u_8[83] = in_8[83] + e1_ext[2][83];
//   assign u_9[83] = in_9[83] + e1_ext[2][83];
//   assign u_1[84] = in_1[84] + e1_ext[0][84];
//   assign u_2[84] = in_2[84] + e1_ext[0][84];
//   assign u_3[84] = in_3[84] + e1_ext[0][84];
//   assign u_4[84] = in_4[84] + e1_ext[1][84];
//   assign u_5[84] = in_5[84] + e1_ext[1][84];
//   assign u_6[84] = in_6[84] + e1_ext[1][84];
//   assign u_7[84] = in_7[84] + e1_ext[2][84];
//   assign u_8[84] = in_8[84] + e1_ext[2][84];
//   assign u_9[84] = in_9[84] + e1_ext[2][84];
//   assign u_1[85] = in_1[85] + e1_ext[0][85];
//   assign u_2[85] = in_2[85] + e1_ext[0][85];
//   assign u_3[85] = in_3[85] + e1_ext[0][85];
//   assign u_4[85] = in_4[85] + e1_ext[1][85];
//   assign u_5[85] = in_5[85] + e1_ext[1][85];
//   assign u_6[85] = in_6[85] + e1_ext[1][85];
//   assign u_7[85] = in_7[85] + e1_ext[2][85];
//   assign u_8[85] = in_8[85] + e1_ext[2][85];
//   assign u_9[85] = in_9[85] + e1_ext[2][85];
//   assign u_1[86] = in_1[86] + e1_ext[0][86];
//   assign u_2[86] = in_2[86] + e1_ext[0][86];
//   assign u_3[86] = in_3[86] + e1_ext[0][86];
//   assign u_4[86] = in_4[86] + e1_ext[1][86];
//   assign u_5[86] = in_5[86] + e1_ext[1][86];
//   assign u_6[86] = in_6[86] + e1_ext[1][86];
//   assign u_7[86] = in_7[86] + e1_ext[2][86];
//   assign u_8[86] = in_8[86] + e1_ext[2][86];
//   assign u_9[86] = in_9[86] + e1_ext[2][86];
//   assign u_1[87] = in_1[87] + e1_ext[0][87];
//   assign u_2[87] = in_2[87] + e1_ext[0][87];
//   assign u_3[87] = in_3[87] + e1_ext[0][87];
//   assign u_4[87] = in_4[87] + e1_ext[1][87];
//   assign u_5[87] = in_5[87] + e1_ext[1][87];
//   assign u_6[87] = in_6[87] + e1_ext[1][87];
//   assign u_7[87] = in_7[87] + e1_ext[2][87];
//   assign u_8[87] = in_8[87] + e1_ext[2][87];
//   assign u_9[87] = in_9[87] + e1_ext[2][87];
//   assign u_1[88] = in_1[88] + e1_ext[0][88];
//   assign u_2[88] = in_2[88] + e1_ext[0][88];
//   assign u_3[88] = in_3[88] + e1_ext[0][88];
//   assign u_4[88] = in_4[88] + e1_ext[1][88];
//   assign u_5[88] = in_5[88] + e1_ext[1][88];
//   assign u_6[88] = in_6[88] + e1_ext[1][88];
//   assign u_7[88] = in_7[88] + e1_ext[2][88];
//   assign u_8[88] = in_8[88] + e1_ext[2][88];
//   assign u_9[88] = in_9[88] + e1_ext[2][88];
//   assign u_1[89] = in_1[89] + e1_ext[0][89];
//   assign u_2[89] = in_2[89] + e1_ext[0][89];
//   assign u_3[89] = in_3[89] + e1_ext[0][89];
//   assign u_4[89] = in_4[89] + e1_ext[1][89];
//   assign u_5[89] = in_5[89] + e1_ext[1][89];
//   assign u_6[89] = in_6[89] + e1_ext[1][89];
//   assign u_7[89] = in_7[89] + e1_ext[2][89];
//   assign u_8[89] = in_8[89] + e1_ext[2][89];
//   assign u_9[89] = in_9[89] + e1_ext[2][89];
//   assign u_1[90] = in_1[90] + e1_ext[0][90];
//   assign u_2[90] = in_2[90] + e1_ext[0][90];
//   assign u_3[90] = in_3[90] + e1_ext[0][90];
//   assign u_4[90] = in_4[90] + e1_ext[1][90];
//   assign u_5[90] = in_5[90] + e1_ext[1][90];
//   assign u_6[90] = in_6[90] + e1_ext[1][90];
//   assign u_7[90] = in_7[90] + e1_ext[2][90];
//   assign u_8[90] = in_8[90] + e1_ext[2][90];
//   assign u_9[90] = in_9[90] + e1_ext[2][90];
//   assign u_1[91] = in_1[91] + e1_ext[0][91];
//   assign u_2[91] = in_2[91] + e1_ext[0][91];
//   assign u_3[91] = in_3[91] + e1_ext[0][91];
//   assign u_4[91] = in_4[91] + e1_ext[1][91];
//   assign u_5[91] = in_5[91] + e1_ext[1][91];
//   assign u_6[91] = in_6[91] + e1_ext[1][91];
//   assign u_7[91] = in_7[91] + e1_ext[2][91];
//   assign u_8[91] = in_8[91] + e1_ext[2][91];
//   assign u_9[91] = in_9[91] + e1_ext[2][91];
//   assign u_1[92] = in_1[92] + e1_ext[0][92];
//   assign u_2[92] = in_2[92] + e1_ext[0][92];
//   assign u_3[92] = in_3[92] + e1_ext[0][92];
//   assign u_4[92] = in_4[92] + e1_ext[1][92];
//   assign u_5[92] = in_5[92] + e1_ext[1][92];
//   assign u_6[92] = in_6[92] + e1_ext[1][92];
//   assign u_7[92] = in_7[92] + e1_ext[2][92];
//   assign u_8[92] = in_8[92] + e1_ext[2][92];
//   assign u_9[92] = in_9[92] + e1_ext[2][92];
//   assign u_1[93] = in_1[93] + e1_ext[0][93];
//   assign u_2[93] = in_2[93] + e1_ext[0][93];
//   assign u_3[93] = in_3[93] + e1_ext[0][93];
//   assign u_4[93] = in_4[93] + e1_ext[1][93];
//   assign u_5[93] = in_5[93] + e1_ext[1][93];
//   assign u_6[93] = in_6[93] + e1_ext[1][93];
//   assign u_7[93] = in_7[93] + e1_ext[2][93];
//   assign u_8[93] = in_8[93] + e1_ext[2][93];
//   assign u_9[93] = in_9[93] + e1_ext[2][93];
//   assign u_1[94] = in_1[94] + e1_ext[0][94];
//   assign u_2[94] = in_2[94] + e1_ext[0][94];
//   assign u_3[94] = in_3[94] + e1_ext[0][94];
//   assign u_4[94] = in_4[94] + e1_ext[1][94];
//   assign u_5[94] = in_5[94] + e1_ext[1][94];
//   assign u_6[94] = in_6[94] + e1_ext[1][94];
//   assign u_7[94] = in_7[94] + e1_ext[2][94];
//   assign u_8[94] = in_8[94] + e1_ext[2][94];
//   assign u_9[94] = in_9[94] + e1_ext[2][94];
//   assign u_1[95] = in_1[95] + e1_ext[0][95];
//   assign u_2[95] = in_2[95] + e1_ext[0][95];
//   assign u_3[95] = in_3[95] + e1_ext[0][95];
//   assign u_4[95] = in_4[95] + e1_ext[1][95];
//   assign u_5[95] = in_5[95] + e1_ext[1][95];
//   assign u_6[95] = in_6[95] + e1_ext[1][95];
//   assign u_7[95] = in_7[95] + e1_ext[2][95];
//   assign u_8[95] = in_8[95] + e1_ext[2][95];
//   assign u_9[95] = in_9[95] + e1_ext[2][95];
//   assign u_1[96] = in_1[96] + e1_ext[0][96];
//   assign u_2[96] = in_2[96] + e1_ext[0][96];
//   assign u_3[96] = in_3[96] + e1_ext[0][96];
//   assign u_4[96] = in_4[96] + e1_ext[1][96];
//   assign u_5[96] = in_5[96] + e1_ext[1][96];
//   assign u_6[96] = in_6[96] + e1_ext[1][96];
//   assign u_7[96] = in_7[96] + e1_ext[2][96];
//   assign u_8[96] = in_8[96] + e1_ext[2][96];
//   assign u_9[96] = in_9[96] + e1_ext[2][96];
//   assign u_1[97] = in_1[97] + e1_ext[0][97];
//   assign u_2[97] = in_2[97] + e1_ext[0][97];
//   assign u_3[97] = in_3[97] + e1_ext[0][97];
//   assign u_4[97] = in_4[97] + e1_ext[1][97];
//   assign u_5[97] = in_5[97] + e1_ext[1][97];
//   assign u_6[97] = in_6[97] + e1_ext[1][97];
//   assign u_7[97] = in_7[97] + e1_ext[2][97];
//   assign u_8[97] = in_8[97] + e1_ext[2][97];
//   assign u_9[97] = in_9[97] + e1_ext[2][97];
//   assign u_1[98] = in_1[98] + e1_ext[0][98];
//   assign u_2[98] = in_2[98] + e1_ext[0][98];
//   assign u_3[98] = in_3[98] + e1_ext[0][98];
//   assign u_4[98] = in_4[98] + e1_ext[1][98];
//   assign u_5[98] = in_5[98] + e1_ext[1][98];
//   assign u_6[98] = in_6[98] + e1_ext[1][98];
//   assign u_7[98] = in_7[98] + e1_ext[2][98];
//   assign u_8[98] = in_8[98] + e1_ext[2][98];
//   assign u_9[98] = in_9[98] + e1_ext[2][98];
//   assign u_1[99] = in_1[99] + e1_ext[0][99];
//   assign u_2[99] = in_2[99] + e1_ext[0][99];
//   assign u_3[99] = in_3[99] + e1_ext[0][99];
//   assign u_4[99] = in_4[99] + e1_ext[1][99];
//   assign u_5[99] = in_5[99] + e1_ext[1][99];
//   assign u_6[99] = in_6[99] + e1_ext[1][99];
//   assign u_7[99] = in_7[99] + e1_ext[2][99];
//   assign u_8[99] = in_8[99] + e1_ext[2][99];
//   assign u_9[99] = in_9[99] + e1_ext[2][99];
//   assign u_1[100] = in_1[100] + e1_ext[0][100];
//   assign u_2[100] = in_2[100] + e1_ext[0][100];
//   assign u_3[100] = in_3[100] + e1_ext[0][100];
//   assign u_4[100] = in_4[100] + e1_ext[1][100];
//   assign u_5[100] = in_5[100] + e1_ext[1][100];
//   assign u_6[100] = in_6[100] + e1_ext[1][100];
//   assign u_7[100] = in_7[100] + e1_ext[2][100];
//   assign u_8[100] = in_8[100] + e1_ext[2][100];
//   assign u_9[100] = in_9[100] + e1_ext[2][100];
//   assign u_1[101] = in_1[101] + e1_ext[0][101];
//   assign u_2[101] = in_2[101] + e1_ext[0][101];
//   assign u_3[101] = in_3[101] + e1_ext[0][101];
//   assign u_4[101] = in_4[101] + e1_ext[1][101];
//   assign u_5[101] = in_5[101] + e1_ext[1][101];
//   assign u_6[101] = in_6[101] + e1_ext[1][101];
//   assign u_7[101] = in_7[101] + e1_ext[2][101];
//   assign u_8[101] = in_8[101] + e1_ext[2][101];
//   assign u_9[101] = in_9[101] + e1_ext[2][101];
//   assign u_1[102] = in_1[102] + e1_ext[0][102];
//   assign u_2[102] = in_2[102] + e1_ext[0][102];
//   assign u_3[102] = in_3[102] + e1_ext[0][102];
//   assign u_4[102] = in_4[102] + e1_ext[1][102];
//   assign u_5[102] = in_5[102] + e1_ext[1][102];
//   assign u_6[102] = in_6[102] + e1_ext[1][102];
//   assign u_7[102] = in_7[102] + e1_ext[2][102];
//   assign u_8[102] = in_8[102] + e1_ext[2][102];
//   assign u_9[102] = in_9[102] + e1_ext[2][102];
//   assign u_1[103] = in_1[103] + e1_ext[0][103];
//   assign u_2[103] = in_2[103] + e1_ext[0][103];
//   assign u_3[103] = in_3[103] + e1_ext[0][103];
//   assign u_4[103] = in_4[103] + e1_ext[1][103];
//   assign u_5[103] = in_5[103] + e1_ext[1][103];
//   assign u_6[103] = in_6[103] + e1_ext[1][103];
//   assign u_7[103] = in_7[103] + e1_ext[2][103];
//   assign u_8[103] = in_8[103] + e1_ext[2][103];
//   assign u_9[103] = in_9[103] + e1_ext[2][103];
//   assign u_1[104] = in_1[104] + e1_ext[0][104];
//   assign u_2[104] = in_2[104] + e1_ext[0][104];
//   assign u_3[104] = in_3[104] + e1_ext[0][104];
//   assign u_4[104] = in_4[104] + e1_ext[1][104];
//   assign u_5[104] = in_5[104] + e1_ext[1][104];
//   assign u_6[104] = in_6[104] + e1_ext[1][104];
//   assign u_7[104] = in_7[104] + e1_ext[2][104];
//   assign u_8[104] = in_8[104] + e1_ext[2][104];
//   assign u_9[104] = in_9[104] + e1_ext[2][104];
//   assign u_1[105] = in_1[105] + e1_ext[0][105];
//   assign u_2[105] = in_2[105] + e1_ext[0][105];
//   assign u_3[105] = in_3[105] + e1_ext[0][105];
//   assign u_4[105] = in_4[105] + e1_ext[1][105];
//   assign u_5[105] = in_5[105] + e1_ext[1][105];
//   assign u_6[105] = in_6[105] + e1_ext[1][105];
//   assign u_7[105] = in_7[105] + e1_ext[2][105];
//   assign u_8[105] = in_8[105] + e1_ext[2][105];
//   assign u_9[105] = in_9[105] + e1_ext[2][105];
//   assign u_1[106] = in_1[106] + e1_ext[0][106];
//   assign u_2[106] = in_2[106] + e1_ext[0][106];
//   assign u_3[106] = in_3[106] + e1_ext[0][106];
//   assign u_4[106] = in_4[106] + e1_ext[1][106];
//   assign u_5[106] = in_5[106] + e1_ext[1][106];
//   assign u_6[106] = in_6[106] + e1_ext[1][106];
//   assign u_7[106] = in_7[106] + e1_ext[2][106];
//   assign u_8[106] = in_8[106] + e1_ext[2][106];
//   assign u_9[106] = in_9[106] + e1_ext[2][106];
//   assign u_1[107] = in_1[107] + e1_ext[0][107];
//   assign u_2[107] = in_2[107] + e1_ext[0][107];
//   assign u_3[107] = in_3[107] + e1_ext[0][107];
//   assign u_4[107] = in_4[107] + e1_ext[1][107];
//   assign u_5[107] = in_5[107] + e1_ext[1][107];
//   assign u_6[107] = in_6[107] + e1_ext[1][107];
//   assign u_7[107] = in_7[107] + e1_ext[2][107];
//   assign u_8[107] = in_8[107] + e1_ext[2][107];
//   assign u_9[107] = in_9[107] + e1_ext[2][107];
//   assign u_1[108] = in_1[108] + e1_ext[0][108];
//   assign u_2[108] = in_2[108] + e1_ext[0][108];
//   assign u_3[108] = in_3[108] + e1_ext[0][108];
//   assign u_4[108] = in_4[108] + e1_ext[1][108];
//   assign u_5[108] = in_5[108] + e1_ext[1][108];
//   assign u_6[108] = in_6[108] + e1_ext[1][108];
//   assign u_7[108] = in_7[108] + e1_ext[2][108];
//   assign u_8[108] = in_8[108] + e1_ext[2][108];
//   assign u_9[108] = in_9[108] + e1_ext[2][108];
//   assign u_1[109] = in_1[109] + e1_ext[0][109];
//   assign u_2[109] = in_2[109] + e1_ext[0][109];
//   assign u_3[109] = in_3[109] + e1_ext[0][109];
//   assign u_4[109] = in_4[109] + e1_ext[1][109];
//   assign u_5[109] = in_5[109] + e1_ext[1][109];
//   assign u_6[109] = in_6[109] + e1_ext[1][109];
//   assign u_7[109] = in_7[109] + e1_ext[2][109];
//   assign u_8[109] = in_8[109] + e1_ext[2][109];
//   assign u_9[109] = in_9[109] + e1_ext[2][109];
//   assign u_1[110] = in_1[110] + e1_ext[0][110];
//   assign u_2[110] = in_2[110] + e1_ext[0][110];
//   assign u_3[110] = in_3[110] + e1_ext[0][110];
//   assign u_4[110] = in_4[110] + e1_ext[1][110];
//   assign u_5[110] = in_5[110] + e1_ext[1][110];
//   assign u_6[110] = in_6[110] + e1_ext[1][110];
//   assign u_7[110] = in_7[110] + e1_ext[2][110];
//   assign u_8[110] = in_8[110] + e1_ext[2][110];
//   assign u_9[110] = in_9[110] + e1_ext[2][110];
//   assign u_1[111] = in_1[111] + e1_ext[0][111];
//   assign u_2[111] = in_2[111] + e1_ext[0][111];
//   assign u_3[111] = in_3[111] + e1_ext[0][111];
//   assign u_4[111] = in_4[111] + e1_ext[1][111];
//   assign u_5[111] = in_5[111] + e1_ext[1][111];
//   assign u_6[111] = in_6[111] + e1_ext[1][111];
//   assign u_7[111] = in_7[111] + e1_ext[2][111];
//   assign u_8[111] = in_8[111] + e1_ext[2][111];
//   assign u_9[111] = in_9[111] + e1_ext[2][111];
//   assign u_1[112] = in_1[112] + e1_ext[0][112];
//   assign u_2[112] = in_2[112] + e1_ext[0][112];
//   assign u_3[112] = in_3[112] + e1_ext[0][112];
//   assign u_4[112] = in_4[112] + e1_ext[1][112];
//   assign u_5[112] = in_5[112] + e1_ext[1][112];
//   assign u_6[112] = in_6[112] + e1_ext[1][112];
//   assign u_7[112] = in_7[112] + e1_ext[2][112];
//   assign u_8[112] = in_8[112] + e1_ext[2][112];
//   assign u_9[112] = in_9[112] + e1_ext[2][112];
//   assign u_1[113] = in_1[113] + e1_ext[0][113];
//   assign u_2[113] = in_2[113] + e1_ext[0][113];
//   assign u_3[113] = in_3[113] + e1_ext[0][113];
//   assign u_4[113] = in_4[113] + e1_ext[1][113];
//   assign u_5[113] = in_5[113] + e1_ext[1][113];
//   assign u_6[113] = in_6[113] + e1_ext[1][113];
//   assign u_7[113] = in_7[113] + e1_ext[2][113];
//   assign u_8[113] = in_8[113] + e1_ext[2][113];
//   assign u_9[113] = in_9[113] + e1_ext[2][113];
//   assign u_1[114] = in_1[114] + e1_ext[0][114];
//   assign u_2[114] = in_2[114] + e1_ext[0][114];
//   assign u_3[114] = in_3[114] + e1_ext[0][114];
//   assign u_4[114] = in_4[114] + e1_ext[1][114];
//   assign u_5[114] = in_5[114] + e1_ext[1][114];
//   assign u_6[114] = in_6[114] + e1_ext[1][114];
//   assign u_7[114] = in_7[114] + e1_ext[2][114];
//   assign u_8[114] = in_8[114] + e1_ext[2][114];
//   assign u_9[114] = in_9[114] + e1_ext[2][114];
//   assign u_1[115] = in_1[115] + e1_ext[0][115];
//   assign u_2[115] = in_2[115] + e1_ext[0][115];
//   assign u_3[115] = in_3[115] + e1_ext[0][115];
//   assign u_4[115] = in_4[115] + e1_ext[1][115];
//   assign u_5[115] = in_5[115] + e1_ext[1][115];
//   assign u_6[115] = in_6[115] + e1_ext[1][115];
//   assign u_7[115] = in_7[115] + e1_ext[2][115];
//   assign u_8[115] = in_8[115] + e1_ext[2][115];
//   assign u_9[115] = in_9[115] + e1_ext[2][115];
//   assign u_1[116] = in_1[116] + e1_ext[0][116];
//   assign u_2[116] = in_2[116] + e1_ext[0][116];
//   assign u_3[116] = in_3[116] + e1_ext[0][116];
//   assign u_4[116] = in_4[116] + e1_ext[1][116];
//   assign u_5[116] = in_5[116] + e1_ext[1][116];
//   assign u_6[116] = in_6[116] + e1_ext[1][116];
//   assign u_7[116] = in_7[116] + e1_ext[2][116];
//   assign u_8[116] = in_8[116] + e1_ext[2][116];
//   assign u_9[116] = in_9[116] + e1_ext[2][116];
//   assign u_1[117] = in_1[117] + e1_ext[0][117];
//   assign u_2[117] = in_2[117] + e1_ext[0][117];
//   assign u_3[117] = in_3[117] + e1_ext[0][117];
//   assign u_4[117] = in_4[117] + e1_ext[1][117];
//   assign u_5[117] = in_5[117] + e1_ext[1][117];
//   assign u_6[117] = in_6[117] + e1_ext[1][117];
//   assign u_7[117] = in_7[117] + e1_ext[2][117];
//   assign u_8[117] = in_8[117] + e1_ext[2][117];
//   assign u_9[117] = in_9[117] + e1_ext[2][117];
//   assign u_1[118] = in_1[118] + e1_ext[0][118];
//   assign u_2[118] = in_2[118] + e1_ext[0][118];
//   assign u_3[118] = in_3[118] + e1_ext[0][118];
//   assign u_4[118] = in_4[118] + e1_ext[1][118];
//   assign u_5[118] = in_5[118] + e1_ext[1][118];
//   assign u_6[118] = in_6[118] + e1_ext[1][118];
//   assign u_7[118] = in_7[118] + e1_ext[2][118];
//   assign u_8[118] = in_8[118] + e1_ext[2][118];
//   assign u_9[118] = in_9[118] + e1_ext[2][118];
//   assign u_1[119] = in_1[119] + e1_ext[0][119];
//   assign u_2[119] = in_2[119] + e1_ext[0][119];
//   assign u_3[119] = in_3[119] + e1_ext[0][119];
//   assign u_4[119] = in_4[119] + e1_ext[1][119];
//   assign u_5[119] = in_5[119] + e1_ext[1][119];
//   assign u_6[119] = in_6[119] + e1_ext[1][119];
//   assign u_7[119] = in_7[119] + e1_ext[2][119];
//   assign u_8[119] = in_8[119] + e1_ext[2][119];
//   assign u_9[119] = in_9[119] + e1_ext[2][119];
//   assign u_1[120] = in_1[120] + e1_ext[0][120];
//   assign u_2[120] = in_2[120] + e1_ext[0][120];
//   assign u_3[120] = in_3[120] + e1_ext[0][120];
//   assign u_4[120] = in_4[120] + e1_ext[1][120];
//   assign u_5[120] = in_5[120] + e1_ext[1][120];
//   assign u_6[120] = in_6[120] + e1_ext[1][120];
//   assign u_7[120] = in_7[120] + e1_ext[2][120];
//   assign u_8[120] = in_8[120] + e1_ext[2][120];
//   assign u_9[120] = in_9[120] + e1_ext[2][120];
//   assign u_1[121] = in_1[121] + e1_ext[0][121];
//   assign u_2[121] = in_2[121] + e1_ext[0][121];
//   assign u_3[121] = in_3[121] + e1_ext[0][121];
//   assign u_4[121] = in_4[121] + e1_ext[1][121];
//   assign u_5[121] = in_5[121] + e1_ext[1][121];
//   assign u_6[121] = in_6[121] + e1_ext[1][121];
//   assign u_7[121] = in_7[121] + e1_ext[2][121];
//   assign u_8[121] = in_8[121] + e1_ext[2][121];
//   assign u_9[121] = in_9[121] + e1_ext[2][121];
//   assign u_1[122] = in_1[122] + e1_ext[0][122];
//   assign u_2[122] = in_2[122] + e1_ext[0][122];
//   assign u_3[122] = in_3[122] + e1_ext[0][122];
//   assign u_4[122] = in_4[122] + e1_ext[1][122];
//   assign u_5[122] = in_5[122] + e1_ext[1][122];
//   assign u_6[122] = in_6[122] + e1_ext[1][122];
//   assign u_7[122] = in_7[122] + e1_ext[2][122];
//   assign u_8[122] = in_8[122] + e1_ext[2][122];
//   assign u_9[122] = in_9[122] + e1_ext[2][122];
//   assign u_1[123] = in_1[123] + e1_ext[0][123];
//   assign u_2[123] = in_2[123] + e1_ext[0][123];
//   assign u_3[123] = in_3[123] + e1_ext[0][123];
//   assign u_4[123] = in_4[123] + e1_ext[1][123];
//   assign u_5[123] = in_5[123] + e1_ext[1][123];
//   assign u_6[123] = in_6[123] + e1_ext[1][123];
//   assign u_7[123] = in_7[123] + e1_ext[2][123];
//   assign u_8[123] = in_8[123] + e1_ext[2][123];
//   assign u_9[123] = in_9[123] + e1_ext[2][123];
//   assign u_1[124] = in_1[124] + e1_ext[0][124];
//   assign u_2[124] = in_2[124] + e1_ext[0][124];
//   assign u_3[124] = in_3[124] + e1_ext[0][124];
//   assign u_4[124] = in_4[124] + e1_ext[1][124];
//   assign u_5[124] = in_5[124] + e1_ext[1][124];
//   assign u_6[124] = in_6[124] + e1_ext[1][124];
//   assign u_7[124] = in_7[124] + e1_ext[2][124];
//   assign u_8[124] = in_8[124] + e1_ext[2][124];
//   assign u_9[124] = in_9[124] + e1_ext[2][124];
//   assign u_1[125] = in_1[125] + e1_ext[0][125];
//   assign u_2[125] = in_2[125] + e1_ext[0][125];
//   assign u_3[125] = in_3[125] + e1_ext[0][125];
//   assign u_4[125] = in_4[125] + e1_ext[1][125];
//   assign u_5[125] = in_5[125] + e1_ext[1][125];
//   assign u_6[125] = in_6[125] + e1_ext[1][125];
//   assign u_7[125] = in_7[125] + e1_ext[2][125];
//   assign u_8[125] = in_8[125] + e1_ext[2][125];
//   assign u_9[125] = in_9[125] + e1_ext[2][125];
//   assign u_1[126] = in_1[126] + e1_ext[0][126];
//   assign u_2[126] = in_2[126] + e1_ext[0][126];
//   assign u_3[126] = in_3[126] + e1_ext[0][126];
//   assign u_4[126] = in_4[126] + e1_ext[1][126];
//   assign u_5[126] = in_5[126] + e1_ext[1][126];
//   assign u_6[126] = in_6[126] + e1_ext[1][126];
//   assign u_7[126] = in_7[126] + e1_ext[2][126];
//   assign u_8[126] = in_8[126] + e1_ext[2][126];
//   assign u_9[126] = in_9[126] + e1_ext[2][126];
//   assign u_1[127] = in_1[127] + e1_ext[0][127];
//   assign u_2[127] = in_2[127] + e1_ext[0][127];
//   assign u_3[127] = in_3[127] + e1_ext[0][127];
//   assign u_4[127] = in_4[127] + e1_ext[1][127];
//   assign u_5[127] = in_5[127] + e1_ext[1][127];
//   assign u_6[127] = in_6[127] + e1_ext[1][127];
//   assign u_7[127] = in_7[127] + e1_ext[2][127];
//   assign u_8[127] = in_8[127] + e1_ext[2][127];
//   assign u_9[127] = in_9[127] + e1_ext[2][127];
//   assign u_1[128] = in_1[128] + e1_ext[0][128];
//   assign u_2[128] = in_2[128] + e1_ext[0][128];
//   assign u_3[128] = in_3[128] + e1_ext[0][128];
//   assign u_4[128] = in_4[128] + e1_ext[1][128];
//   assign u_5[128] = in_5[128] + e1_ext[1][128];
//   assign u_6[128] = in_6[128] + e1_ext[1][128];
//   assign u_7[128] = in_7[128] + e1_ext[2][128];
//   assign u_8[128] = in_8[128] + e1_ext[2][128];
//   assign u_9[128] = in_9[128] + e1_ext[2][128];
//   assign u_1[129] = in_1[129] + e1_ext[0][129];
//   assign u_2[129] = in_2[129] + e1_ext[0][129];
//   assign u_3[129] = in_3[129] + e1_ext[0][129];
//   assign u_4[129] = in_4[129] + e1_ext[1][129];
//   assign u_5[129] = in_5[129] + e1_ext[1][129];
//   assign u_6[129] = in_6[129] + e1_ext[1][129];
//   assign u_7[129] = in_7[129] + e1_ext[2][129];
//   assign u_8[129] = in_8[129] + e1_ext[2][129];
//   assign u_9[129] = in_9[129] + e1_ext[2][129];
//   assign u_1[130] = in_1[130] + e1_ext[0][130];
//   assign u_2[130] = in_2[130] + e1_ext[0][130];
//   assign u_3[130] = in_3[130] + e1_ext[0][130];
//   assign u_4[130] = in_4[130] + e1_ext[1][130];
//   assign u_5[130] = in_5[130] + e1_ext[1][130];
//   assign u_6[130] = in_6[130] + e1_ext[1][130];
//   assign u_7[130] = in_7[130] + e1_ext[2][130];
//   assign u_8[130] = in_8[130] + e1_ext[2][130];
//   assign u_9[130] = in_9[130] + e1_ext[2][130];
//   assign u_1[131] = in_1[131] + e1_ext[0][131];
//   assign u_2[131] = in_2[131] + e1_ext[0][131];
//   assign u_3[131] = in_3[131] + e1_ext[0][131];
//   assign u_4[131] = in_4[131] + e1_ext[1][131];
//   assign u_5[131] = in_5[131] + e1_ext[1][131];
//   assign u_6[131] = in_6[131] + e1_ext[1][131];
//   assign u_7[131] = in_7[131] + e1_ext[2][131];
//   assign u_8[131] = in_8[131] + e1_ext[2][131];
//   assign u_9[131] = in_9[131] + e1_ext[2][131];
//   assign u_1[132] = in_1[132] + e1_ext[0][132];
//   assign u_2[132] = in_2[132] + e1_ext[0][132];
//   assign u_3[132] = in_3[132] + e1_ext[0][132];
//   assign u_4[132] = in_4[132] + e1_ext[1][132];
//   assign u_5[132] = in_5[132] + e1_ext[1][132];
//   assign u_6[132] = in_6[132] + e1_ext[1][132];
//   assign u_7[132] = in_7[132] + e1_ext[2][132];
//   assign u_8[132] = in_8[132] + e1_ext[2][132];
//   assign u_9[132] = in_9[132] + e1_ext[2][132];
//   assign u_1[133] = in_1[133] + e1_ext[0][133];
//   assign u_2[133] = in_2[133] + e1_ext[0][133];
//   assign u_3[133] = in_3[133] + e1_ext[0][133];
//   assign u_4[133] = in_4[133] + e1_ext[1][133];
//   assign u_5[133] = in_5[133] + e1_ext[1][133];
//   assign u_6[133] = in_6[133] + e1_ext[1][133];
//   assign u_7[133] = in_7[133] + e1_ext[2][133];
//   assign u_8[133] = in_8[133] + e1_ext[2][133];
//   assign u_9[133] = in_9[133] + e1_ext[2][133];
//   assign u_1[134] = in_1[134] + e1_ext[0][134];
//   assign u_2[134] = in_2[134] + e1_ext[0][134];
//   assign u_3[134] = in_3[134] + e1_ext[0][134];
//   assign u_4[134] = in_4[134] + e1_ext[1][134];
//   assign u_5[134] = in_5[134] + e1_ext[1][134];
//   assign u_6[134] = in_6[134] + e1_ext[1][134];
//   assign u_7[134] = in_7[134] + e1_ext[2][134];
//   assign u_8[134] = in_8[134] + e1_ext[2][134];
//   assign u_9[134] = in_9[134] + e1_ext[2][134];
//   assign u_1[135] = in_1[135] + e1_ext[0][135];
//   assign u_2[135] = in_2[135] + e1_ext[0][135];
//   assign u_3[135] = in_3[135] + e1_ext[0][135];
//   assign u_4[135] = in_4[135] + e1_ext[1][135];
//   assign u_5[135] = in_5[135] + e1_ext[1][135];
//   assign u_6[135] = in_6[135] + e1_ext[1][135];
//   assign u_7[135] = in_7[135] + e1_ext[2][135];
//   assign u_8[135] = in_8[135] + e1_ext[2][135];
//   assign u_9[135] = in_9[135] + e1_ext[2][135];
//   assign u_1[136] = in_1[136] + e1_ext[0][136];
//   assign u_2[136] = in_2[136] + e1_ext[0][136];
//   assign u_3[136] = in_3[136] + e1_ext[0][136];
//   assign u_4[136] = in_4[136] + e1_ext[1][136];
//   assign u_5[136] = in_5[136] + e1_ext[1][136];
//   assign u_6[136] = in_6[136] + e1_ext[1][136];
//   assign u_7[136] = in_7[136] + e1_ext[2][136];
//   assign u_8[136] = in_8[136] + e1_ext[2][136];
//   assign u_9[136] = in_9[136] + e1_ext[2][136];
//   assign u_1[137] = in_1[137] + e1_ext[0][137];
//   assign u_2[137] = in_2[137] + e1_ext[0][137];
//   assign u_3[137] = in_3[137] + e1_ext[0][137];
//   assign u_4[137] = in_4[137] + e1_ext[1][137];
//   assign u_5[137] = in_5[137] + e1_ext[1][137];
//   assign u_6[137] = in_6[137] + e1_ext[1][137];
//   assign u_7[137] = in_7[137] + e1_ext[2][137];
//   assign u_8[137] = in_8[137] + e1_ext[2][137];
//   assign u_9[137] = in_9[137] + e1_ext[2][137];
//   assign u_1[138] = in_1[138] + e1_ext[0][138];
//   assign u_2[138] = in_2[138] + e1_ext[0][138];
//   assign u_3[138] = in_3[138] + e1_ext[0][138];
//   assign u_4[138] = in_4[138] + e1_ext[1][138];
//   assign u_5[138] = in_5[138] + e1_ext[1][138];
//   assign u_6[138] = in_6[138] + e1_ext[1][138];
//   assign u_7[138] = in_7[138] + e1_ext[2][138];
//   assign u_8[138] = in_8[138] + e1_ext[2][138];
//   assign u_9[138] = in_9[138] + e1_ext[2][138];
//   assign u_1[139] = in_1[139] + e1_ext[0][139];
//   assign u_2[139] = in_2[139] + e1_ext[0][139];
//   assign u_3[139] = in_3[139] + e1_ext[0][139];
//   assign u_4[139] = in_4[139] + e1_ext[1][139];
//   assign u_5[139] = in_5[139] + e1_ext[1][139];
//   assign u_6[139] = in_6[139] + e1_ext[1][139];
//   assign u_7[139] = in_7[139] + e1_ext[2][139];
//   assign u_8[139] = in_8[139] + e1_ext[2][139];
//   assign u_9[139] = in_9[139] + e1_ext[2][139];
//   assign u_1[140] = in_1[140] + e1_ext[0][140];
//   assign u_2[140] = in_2[140] + e1_ext[0][140];
//   assign u_3[140] = in_3[140] + e1_ext[0][140];
//   assign u_4[140] = in_4[140] + e1_ext[1][140];
//   assign u_5[140] = in_5[140] + e1_ext[1][140];
//   assign u_6[140] = in_6[140] + e1_ext[1][140];
//   assign u_7[140] = in_7[140] + e1_ext[2][140];
//   assign u_8[140] = in_8[140] + e1_ext[2][140];
//   assign u_9[140] = in_9[140] + e1_ext[2][140];
//   assign u_1[141] = in_1[141] + e1_ext[0][141];
//   assign u_2[141] = in_2[141] + e1_ext[0][141];
//   assign u_3[141] = in_3[141] + e1_ext[0][141];
//   assign u_4[141] = in_4[141] + e1_ext[1][141];
//   assign u_5[141] = in_5[141] + e1_ext[1][141];
//   assign u_6[141] = in_6[141] + e1_ext[1][141];
//   assign u_7[141] = in_7[141] + e1_ext[2][141];
//   assign u_8[141] = in_8[141] + e1_ext[2][141];
//   assign u_9[141] = in_9[141] + e1_ext[2][141];
//   assign u_1[142] = in_1[142] + e1_ext[0][142];
//   assign u_2[142] = in_2[142] + e1_ext[0][142];
//   assign u_3[142] = in_3[142] + e1_ext[0][142];
//   assign u_4[142] = in_4[142] + e1_ext[1][142];
//   assign u_5[142] = in_5[142] + e1_ext[1][142];
//   assign u_6[142] = in_6[142] + e1_ext[1][142];
//   assign u_7[142] = in_7[142] + e1_ext[2][142];
//   assign u_8[142] = in_8[142] + e1_ext[2][142];
//   assign u_9[142] = in_9[142] + e1_ext[2][142];
//   assign u_1[143] = in_1[143] + e1_ext[0][143];
//   assign u_2[143] = in_2[143] + e1_ext[0][143];
//   assign u_3[143] = in_3[143] + e1_ext[0][143];
//   assign u_4[143] = in_4[143] + e1_ext[1][143];
//   assign u_5[143] = in_5[143] + e1_ext[1][143];
//   assign u_6[143] = in_6[143] + e1_ext[1][143];
//   assign u_7[143] = in_7[143] + e1_ext[2][143];
//   assign u_8[143] = in_8[143] + e1_ext[2][143];
//   assign u_9[143] = in_9[143] + e1_ext[2][143];
//   assign u_1[144] = in_1[144] + e1_ext[0][144];
//   assign u_2[144] = in_2[144] + e1_ext[0][144];
//   assign u_3[144] = in_3[144] + e1_ext[0][144];
//   assign u_4[144] = in_4[144] + e1_ext[1][144];
//   assign u_5[144] = in_5[144] + e1_ext[1][144];
//   assign u_6[144] = in_6[144] + e1_ext[1][144];
//   assign u_7[144] = in_7[144] + e1_ext[2][144];
//   assign u_8[144] = in_8[144] + e1_ext[2][144];
//   assign u_9[144] = in_9[144] + e1_ext[2][144];
//   assign u_1[145] = in_1[145] + e1_ext[0][145];
//   assign u_2[145] = in_2[145] + e1_ext[0][145];
//   assign u_3[145] = in_3[145] + e1_ext[0][145];
//   assign u_4[145] = in_4[145] + e1_ext[1][145];
//   assign u_5[145] = in_5[145] + e1_ext[1][145];
//   assign u_6[145] = in_6[145] + e1_ext[1][145];
//   assign u_7[145] = in_7[145] + e1_ext[2][145];
//   assign u_8[145] = in_8[145] + e1_ext[2][145];
//   assign u_9[145] = in_9[145] + e1_ext[2][145];
//   assign u_1[146] = in_1[146] + e1_ext[0][146];
//   assign u_2[146] = in_2[146] + e1_ext[0][146];
//   assign u_3[146] = in_3[146] + e1_ext[0][146];
//   assign u_4[146] = in_4[146] + e1_ext[1][146];
//   assign u_5[146] = in_5[146] + e1_ext[1][146];
//   assign u_6[146] = in_6[146] + e1_ext[1][146];
//   assign u_7[146] = in_7[146] + e1_ext[2][146];
//   assign u_8[146] = in_8[146] + e1_ext[2][146];
//   assign u_9[146] = in_9[146] + e1_ext[2][146];
//   assign u_1[147] = in_1[147] + e1_ext[0][147];
//   assign u_2[147] = in_2[147] + e1_ext[0][147];
//   assign u_3[147] = in_3[147] + e1_ext[0][147];
//   assign u_4[147] = in_4[147] + e1_ext[1][147];
//   assign u_5[147] = in_5[147] + e1_ext[1][147];
//   assign u_6[147] = in_6[147] + e1_ext[1][147];
//   assign u_7[147] = in_7[147] + e1_ext[2][147];
//   assign u_8[147] = in_8[147] + e1_ext[2][147];
//   assign u_9[147] = in_9[147] + e1_ext[2][147];
//   assign u_1[148] = in_1[148] + e1_ext[0][148];
//   assign u_2[148] = in_2[148] + e1_ext[0][148];
//   assign u_3[148] = in_3[148] + e1_ext[0][148];
//   assign u_4[148] = in_4[148] + e1_ext[1][148];
//   assign u_5[148] = in_5[148] + e1_ext[1][148];
//   assign u_6[148] = in_6[148] + e1_ext[1][148];
//   assign u_7[148] = in_7[148] + e1_ext[2][148];
//   assign u_8[148] = in_8[148] + e1_ext[2][148];
//   assign u_9[148] = in_9[148] + e1_ext[2][148];
//   assign u_1[149] = in_1[149] + e1_ext[0][149];
//   assign u_2[149] = in_2[149] + e1_ext[0][149];
//   assign u_3[149] = in_3[149] + e1_ext[0][149];
//   assign u_4[149] = in_4[149] + e1_ext[1][149];
//   assign u_5[149] = in_5[149] + e1_ext[1][149];
//   assign u_6[149] = in_6[149] + e1_ext[1][149];
//   assign u_7[149] = in_7[149] + e1_ext[2][149];
//   assign u_8[149] = in_8[149] + e1_ext[2][149];
//   assign u_9[149] = in_9[149] + e1_ext[2][149];
//   assign u_1[150] = in_1[150] + e1_ext[0][150];
//   assign u_2[150] = in_2[150] + e1_ext[0][150];
//   assign u_3[150] = in_3[150] + e1_ext[0][150];
//   assign u_4[150] = in_4[150] + e1_ext[1][150];
//   assign u_5[150] = in_5[150] + e1_ext[1][150];
//   assign u_6[150] = in_6[150] + e1_ext[1][150];
//   assign u_7[150] = in_7[150] + e1_ext[2][150];
//   assign u_8[150] = in_8[150] + e1_ext[2][150];
//   assign u_9[150] = in_9[150] + e1_ext[2][150];
//   assign u_1[151] = in_1[151] + e1_ext[0][151];
//   assign u_2[151] = in_2[151] + e1_ext[0][151];
//   assign u_3[151] = in_3[151] + e1_ext[0][151];
//   assign u_4[151] = in_4[151] + e1_ext[1][151];
//   assign u_5[151] = in_5[151] + e1_ext[1][151];
//   assign u_6[151] = in_6[151] + e1_ext[1][151];
//   assign u_7[151] = in_7[151] + e1_ext[2][151];
//   assign u_8[151] = in_8[151] + e1_ext[2][151];
//   assign u_9[151] = in_9[151] + e1_ext[2][151];
//   assign u_1[152] = in_1[152] + e1_ext[0][152];
//   assign u_2[152] = in_2[152] + e1_ext[0][152];
//   assign u_3[152] = in_3[152] + e1_ext[0][152];
//   assign u_4[152] = in_4[152] + e1_ext[1][152];
//   assign u_5[152] = in_5[152] + e1_ext[1][152];
//   assign u_6[152] = in_6[152] + e1_ext[1][152];
//   assign u_7[152] = in_7[152] + e1_ext[2][152];
//   assign u_8[152] = in_8[152] + e1_ext[2][152];
//   assign u_9[152] = in_9[152] + e1_ext[2][152];
//   assign u_1[153] = in_1[153] + e1_ext[0][153];
//   assign u_2[153] = in_2[153] + e1_ext[0][153];
//   assign u_3[153] = in_3[153] + e1_ext[0][153];
//   assign u_4[153] = in_4[153] + e1_ext[1][153];
//   assign u_5[153] = in_5[153] + e1_ext[1][153];
//   assign u_6[153] = in_6[153] + e1_ext[1][153];
//   assign u_7[153] = in_7[153] + e1_ext[2][153];
//   assign u_8[153] = in_8[153] + e1_ext[2][153];
//   assign u_9[153] = in_9[153] + e1_ext[2][153];
//   assign u_1[154] = in_1[154] + e1_ext[0][154];
//   assign u_2[154] = in_2[154] + e1_ext[0][154];
//   assign u_3[154] = in_3[154] + e1_ext[0][154];
//   assign u_4[154] = in_4[154] + e1_ext[1][154];
//   assign u_5[154] = in_5[154] + e1_ext[1][154];
//   assign u_6[154] = in_6[154] + e1_ext[1][154];
//   assign u_7[154] = in_7[154] + e1_ext[2][154];
//   assign u_8[154] = in_8[154] + e1_ext[2][154];
//   assign u_9[154] = in_9[154] + e1_ext[2][154];
//   assign u_1[155] = in_1[155] + e1_ext[0][155];
//   assign u_2[155] = in_2[155] + e1_ext[0][155];
//   assign u_3[155] = in_3[155] + e1_ext[0][155];
//   assign u_4[155] = in_4[155] + e1_ext[1][155];
//   assign u_5[155] = in_5[155] + e1_ext[1][155];
//   assign u_6[155] = in_6[155] + e1_ext[1][155];
//   assign u_7[155] = in_7[155] + e1_ext[2][155];
//   assign u_8[155] = in_8[155] + e1_ext[2][155];
//   assign u_9[155] = in_9[155] + e1_ext[2][155];
//   assign u_1[156] = in_1[156] + e1_ext[0][156];
//   assign u_2[156] = in_2[156] + e1_ext[0][156];
//   assign u_3[156] = in_3[156] + e1_ext[0][156];
//   assign u_4[156] = in_4[156] + e1_ext[1][156];
//   assign u_5[156] = in_5[156] + e1_ext[1][156];
//   assign u_6[156] = in_6[156] + e1_ext[1][156];
//   assign u_7[156] = in_7[156] + e1_ext[2][156];
//   assign u_8[156] = in_8[156] + e1_ext[2][156];
//   assign u_9[156] = in_9[156] + e1_ext[2][156];
//   assign u_1[157] = in_1[157] + e1_ext[0][157];
//   assign u_2[157] = in_2[157] + e1_ext[0][157];
//   assign u_3[157] = in_3[157] + e1_ext[0][157];
//   assign u_4[157] = in_4[157] + e1_ext[1][157];
//   assign u_5[157] = in_5[157] + e1_ext[1][157];
//   assign u_6[157] = in_6[157] + e1_ext[1][157];
//   assign u_7[157] = in_7[157] + e1_ext[2][157];
//   assign u_8[157] = in_8[157] + e1_ext[2][157];
//   assign u_9[157] = in_9[157] + e1_ext[2][157];
//   assign u_1[158] = in_1[158] + e1_ext[0][158];
//   assign u_2[158] = in_2[158] + e1_ext[0][158];
//   assign u_3[158] = in_3[158] + e1_ext[0][158];
//   assign u_4[158] = in_4[158] + e1_ext[1][158];
//   assign u_5[158] = in_5[158] + e1_ext[1][158];
//   assign u_6[158] = in_6[158] + e1_ext[1][158];
//   assign u_7[158] = in_7[158] + e1_ext[2][158];
//   assign u_8[158] = in_8[158] + e1_ext[2][158];
//   assign u_9[158] = in_9[158] + e1_ext[2][158];
//   assign u_1[159] = in_1[159] + e1_ext[0][159];
//   assign u_2[159] = in_2[159] + e1_ext[0][159];
//   assign u_3[159] = in_3[159] + e1_ext[0][159];
//   assign u_4[159] = in_4[159] + e1_ext[1][159];
//   assign u_5[159] = in_5[159] + e1_ext[1][159];
//   assign u_6[159] = in_6[159] + e1_ext[1][159];
//   assign u_7[159] = in_7[159] + e1_ext[2][159];
//   assign u_8[159] = in_8[159] + e1_ext[2][159];
//   assign u_9[159] = in_9[159] + e1_ext[2][159];
//   assign u_1[160] = in_1[160] + e1_ext[0][160];
//   assign u_2[160] = in_2[160] + e1_ext[0][160];
//   assign u_3[160] = in_3[160] + e1_ext[0][160];
//   assign u_4[160] = in_4[160] + e1_ext[1][160];
//   assign u_5[160] = in_5[160] + e1_ext[1][160];
//   assign u_6[160] = in_6[160] + e1_ext[1][160];
//   assign u_7[160] = in_7[160] + e1_ext[2][160];
//   assign u_8[160] = in_8[160] + e1_ext[2][160];
//   assign u_9[160] = in_9[160] + e1_ext[2][160];
//   assign u_1[161] = in_1[161] + e1_ext[0][161];
//   assign u_2[161] = in_2[161] + e1_ext[0][161];
//   assign u_3[161] = in_3[161] + e1_ext[0][161];
//   assign u_4[161] = in_4[161] + e1_ext[1][161];
//   assign u_5[161] = in_5[161] + e1_ext[1][161];
//   assign u_6[161] = in_6[161] + e1_ext[1][161];
//   assign u_7[161] = in_7[161] + e1_ext[2][161];
//   assign u_8[161] = in_8[161] + e1_ext[2][161];
//   assign u_9[161] = in_9[161] + e1_ext[2][161];
//   assign u_1[162] = in_1[162] + e1_ext[0][162];
//   assign u_2[162] = in_2[162] + e1_ext[0][162];
//   assign u_3[162] = in_3[162] + e1_ext[0][162];
//   assign u_4[162] = in_4[162] + e1_ext[1][162];
//   assign u_5[162] = in_5[162] + e1_ext[1][162];
//   assign u_6[162] = in_6[162] + e1_ext[1][162];
//   assign u_7[162] = in_7[162] + e1_ext[2][162];
//   assign u_8[162] = in_8[162] + e1_ext[2][162];
//   assign u_9[162] = in_9[162] + e1_ext[2][162];
//   assign u_1[163] = in_1[163] + e1_ext[0][163];
//   assign u_2[163] = in_2[163] + e1_ext[0][163];
//   assign u_3[163] = in_3[163] + e1_ext[0][163];
//   assign u_4[163] = in_4[163] + e1_ext[1][163];
//   assign u_5[163] = in_5[163] + e1_ext[1][163];
//   assign u_6[163] = in_6[163] + e1_ext[1][163];
//   assign u_7[163] = in_7[163] + e1_ext[2][163];
//   assign u_8[163] = in_8[163] + e1_ext[2][163];
//   assign u_9[163] = in_9[163] + e1_ext[2][163];
//   assign u_1[164] = in_1[164] + e1_ext[0][164];
//   assign u_2[164] = in_2[164] + e1_ext[0][164];
//   assign u_3[164] = in_3[164] + e1_ext[0][164];
//   assign u_4[164] = in_4[164] + e1_ext[1][164];
//   assign u_5[164] = in_5[164] + e1_ext[1][164];
//   assign u_6[164] = in_6[164] + e1_ext[1][164];
//   assign u_7[164] = in_7[164] + e1_ext[2][164];
//   assign u_8[164] = in_8[164] + e1_ext[2][164];
//   assign u_9[164] = in_9[164] + e1_ext[2][164];
//   assign u_1[165] = in_1[165] + e1_ext[0][165];
//   assign u_2[165] = in_2[165] + e1_ext[0][165];
//   assign u_3[165] = in_3[165] + e1_ext[0][165];
//   assign u_4[165] = in_4[165] + e1_ext[1][165];
//   assign u_5[165] = in_5[165] + e1_ext[1][165];
//   assign u_6[165] = in_6[165] + e1_ext[1][165];
//   assign u_7[165] = in_7[165] + e1_ext[2][165];
//   assign u_8[165] = in_8[165] + e1_ext[2][165];
//   assign u_9[165] = in_9[165] + e1_ext[2][165];
//   assign u_1[166] = in_1[166] + e1_ext[0][166];
//   assign u_2[166] = in_2[166] + e1_ext[0][166];
//   assign u_3[166] = in_3[166] + e1_ext[0][166];
//   assign u_4[166] = in_4[166] + e1_ext[1][166];
//   assign u_5[166] = in_5[166] + e1_ext[1][166];
//   assign u_6[166] = in_6[166] + e1_ext[1][166];
//   assign u_7[166] = in_7[166] + e1_ext[2][166];
//   assign u_8[166] = in_8[166] + e1_ext[2][166];
//   assign u_9[166] = in_9[166] + e1_ext[2][166];
//   assign u_1[167] = in_1[167] + e1_ext[0][167];
//   assign u_2[167] = in_2[167] + e1_ext[0][167];
//   assign u_3[167] = in_3[167] + e1_ext[0][167];
//   assign u_4[167] = in_4[167] + e1_ext[1][167];
//   assign u_5[167] = in_5[167] + e1_ext[1][167];
//   assign u_6[167] = in_6[167] + e1_ext[1][167];
//   assign u_7[167] = in_7[167] + e1_ext[2][167];
//   assign u_8[167] = in_8[167] + e1_ext[2][167];
//   assign u_9[167] = in_9[167] + e1_ext[2][167];
//   assign u_1[168] = in_1[168] + e1_ext[0][168];
//   assign u_2[168] = in_2[168] + e1_ext[0][168];
//   assign u_3[168] = in_3[168] + e1_ext[0][168];
//   assign u_4[168] = in_4[168] + e1_ext[1][168];
//   assign u_5[168] = in_5[168] + e1_ext[1][168];
//   assign u_6[168] = in_6[168] + e1_ext[1][168];
//   assign u_7[168] = in_7[168] + e1_ext[2][168];
//   assign u_8[168] = in_8[168] + e1_ext[2][168];
//   assign u_9[168] = in_9[168] + e1_ext[2][168];
//   assign u_1[169] = in_1[169] + e1_ext[0][169];
//   assign u_2[169] = in_2[169] + e1_ext[0][169];
//   assign u_3[169] = in_3[169] + e1_ext[0][169];
//   assign u_4[169] = in_4[169] + e1_ext[1][169];
//   assign u_5[169] = in_5[169] + e1_ext[1][169];
//   assign u_6[169] = in_6[169] + e1_ext[1][169];
//   assign u_7[169] = in_7[169] + e1_ext[2][169];
//   assign u_8[169] = in_8[169] + e1_ext[2][169];
//   assign u_9[169] = in_9[169] + e1_ext[2][169];
//   assign u_1[170] = in_1[170] + e1_ext[0][170];
//   assign u_2[170] = in_2[170] + e1_ext[0][170];
//   assign u_3[170] = in_3[170] + e1_ext[0][170];
//   assign u_4[170] = in_4[170] + e1_ext[1][170];
//   assign u_5[170] = in_5[170] + e1_ext[1][170];
//   assign u_6[170] = in_6[170] + e1_ext[1][170];
//   assign u_7[170] = in_7[170] + e1_ext[2][170];
//   assign u_8[170] = in_8[170] + e1_ext[2][170];
//   assign u_9[170] = in_9[170] + e1_ext[2][170];
//   assign u_1[171] = in_1[171] + e1_ext[0][171];
//   assign u_2[171] = in_2[171] + e1_ext[0][171];
//   assign u_3[171] = in_3[171] + e1_ext[0][171];
//   assign u_4[171] = in_4[171] + e1_ext[1][171];
//   assign u_5[171] = in_5[171] + e1_ext[1][171];
//   assign u_6[171] = in_6[171] + e1_ext[1][171];
//   assign u_7[171] = in_7[171] + e1_ext[2][171];
//   assign u_8[171] = in_8[171] + e1_ext[2][171];
//   assign u_9[171] = in_9[171] + e1_ext[2][171];
//   assign u_1[172] = in_1[172] + e1_ext[0][172];
//   assign u_2[172] = in_2[172] + e1_ext[0][172];
//   assign u_3[172] = in_3[172] + e1_ext[0][172];
//   assign u_4[172] = in_4[172] + e1_ext[1][172];
//   assign u_5[172] = in_5[172] + e1_ext[1][172];
//   assign u_6[172] = in_6[172] + e1_ext[1][172];
//   assign u_7[172] = in_7[172] + e1_ext[2][172];
//   assign u_8[172] = in_8[172] + e1_ext[2][172];
//   assign u_9[172] = in_9[172] + e1_ext[2][172];
//   assign u_1[173] = in_1[173] + e1_ext[0][173];
//   assign u_2[173] = in_2[173] + e1_ext[0][173];
//   assign u_3[173] = in_3[173] + e1_ext[0][173];
//   assign u_4[173] = in_4[173] + e1_ext[1][173];
//   assign u_5[173] = in_5[173] + e1_ext[1][173];
//   assign u_6[173] = in_6[173] + e1_ext[1][173];
//   assign u_7[173] = in_7[173] + e1_ext[2][173];
//   assign u_8[173] = in_8[173] + e1_ext[2][173];
//   assign u_9[173] = in_9[173] + e1_ext[2][173];
//   assign u_1[174] = in_1[174] + e1_ext[0][174];
//   assign u_2[174] = in_2[174] + e1_ext[0][174];
//   assign u_3[174] = in_3[174] + e1_ext[0][174];
//   assign u_4[174] = in_4[174] + e1_ext[1][174];
//   assign u_5[174] = in_5[174] + e1_ext[1][174];
//   assign u_6[174] = in_6[174] + e1_ext[1][174];
//   assign u_7[174] = in_7[174] + e1_ext[2][174];
//   assign u_8[174] = in_8[174] + e1_ext[2][174];
//   assign u_9[174] = in_9[174] + e1_ext[2][174];
//   assign u_1[175] = in_1[175] + e1_ext[0][175];
//   assign u_2[175] = in_2[175] + e1_ext[0][175];
//   assign u_3[175] = in_3[175] + e1_ext[0][175];
//   assign u_4[175] = in_4[175] + e1_ext[1][175];
//   assign u_5[175] = in_5[175] + e1_ext[1][175];
//   assign u_6[175] = in_6[175] + e1_ext[1][175];
//   assign u_7[175] = in_7[175] + e1_ext[2][175];
//   assign u_8[175] = in_8[175] + e1_ext[2][175];
//   assign u_9[175] = in_9[175] + e1_ext[2][175];
//   assign u_1[176] = in_1[176] + e1_ext[0][176];
//   assign u_2[176] = in_2[176] + e1_ext[0][176];
//   assign u_3[176] = in_3[176] + e1_ext[0][176];
//   assign u_4[176] = in_4[176] + e1_ext[1][176];
//   assign u_5[176] = in_5[176] + e1_ext[1][176];
//   assign u_6[176] = in_6[176] + e1_ext[1][176];
//   assign u_7[176] = in_7[176] + e1_ext[2][176];
//   assign u_8[176] = in_8[176] + e1_ext[2][176];
//   assign u_9[176] = in_9[176] + e1_ext[2][176];
//   assign u_1[177] = in_1[177] + e1_ext[0][177];
//   assign u_2[177] = in_2[177] + e1_ext[0][177];
//   assign u_3[177] = in_3[177] + e1_ext[0][177];
//   assign u_4[177] = in_4[177] + e1_ext[1][177];
//   assign u_5[177] = in_5[177] + e1_ext[1][177];
//   assign u_6[177] = in_6[177] + e1_ext[1][177];
//   assign u_7[177] = in_7[177] + e1_ext[2][177];
//   assign u_8[177] = in_8[177] + e1_ext[2][177];
//   assign u_9[177] = in_9[177] + e1_ext[2][177];
//   assign u_1[178] = in_1[178] + e1_ext[0][178];
//   assign u_2[178] = in_2[178] + e1_ext[0][178];
//   assign u_3[178] = in_3[178] + e1_ext[0][178];
//   assign u_4[178] = in_4[178] + e1_ext[1][178];
//   assign u_5[178] = in_5[178] + e1_ext[1][178];
//   assign u_6[178] = in_6[178] + e1_ext[1][178];
//   assign u_7[178] = in_7[178] + e1_ext[2][178];
//   assign u_8[178] = in_8[178] + e1_ext[2][178];
//   assign u_9[178] = in_9[178] + e1_ext[2][178];
//   assign u_1[179] = in_1[179] + e1_ext[0][179];
//   assign u_2[179] = in_2[179] + e1_ext[0][179];
//   assign u_3[179] = in_3[179] + e1_ext[0][179];
//   assign u_4[179] = in_4[179] + e1_ext[1][179];
//   assign u_5[179] = in_5[179] + e1_ext[1][179];
//   assign u_6[179] = in_6[179] + e1_ext[1][179];
//   assign u_7[179] = in_7[179] + e1_ext[2][179];
//   assign u_8[179] = in_8[179] + e1_ext[2][179];
//   assign u_9[179] = in_9[179] + e1_ext[2][179];
//   assign u_1[180] = in_1[180] + e1_ext[0][180];
//   assign u_2[180] = in_2[180] + e1_ext[0][180];
//   assign u_3[180] = in_3[180] + e1_ext[0][180];
//   assign u_4[180] = in_4[180] + e1_ext[1][180];
//   assign u_5[180] = in_5[180] + e1_ext[1][180];
//   assign u_6[180] = in_6[180] + e1_ext[1][180];
//   assign u_7[180] = in_7[180] + e1_ext[2][180];
//   assign u_8[180] = in_8[180] + e1_ext[2][180];
//   assign u_9[180] = in_9[180] + e1_ext[2][180];
//   assign u_1[181] = in_1[181] + e1_ext[0][181];
//   assign u_2[181] = in_2[181] + e1_ext[0][181];
//   assign u_3[181] = in_3[181] + e1_ext[0][181];
//   assign u_4[181] = in_4[181] + e1_ext[1][181];
//   assign u_5[181] = in_5[181] + e1_ext[1][181];
//   assign u_6[181] = in_6[181] + e1_ext[1][181];
//   assign u_7[181] = in_7[181] + e1_ext[2][181];
//   assign u_8[181] = in_8[181] + e1_ext[2][181];
//   assign u_9[181] = in_9[181] + e1_ext[2][181];
//   assign u_1[182] = in_1[182] + e1_ext[0][182];
//   assign u_2[182] = in_2[182] + e1_ext[0][182];
//   assign u_3[182] = in_3[182] + e1_ext[0][182];
//   assign u_4[182] = in_4[182] + e1_ext[1][182];
//   assign u_5[182] = in_5[182] + e1_ext[1][182];
//   assign u_6[182] = in_6[182] + e1_ext[1][182];
//   assign u_7[182] = in_7[182] + e1_ext[2][182];
//   assign u_8[182] = in_8[182] + e1_ext[2][182];
//   assign u_9[182] = in_9[182] + e1_ext[2][182];
//   assign u_1[183] = in_1[183] + e1_ext[0][183];
//   assign u_2[183] = in_2[183] + e1_ext[0][183];
//   assign u_3[183] = in_3[183] + e1_ext[0][183];
//   assign u_4[183] = in_4[183] + e1_ext[1][183];
//   assign u_5[183] = in_5[183] + e1_ext[1][183];
//   assign u_6[183] = in_6[183] + e1_ext[1][183];
//   assign u_7[183] = in_7[183] + e1_ext[2][183];
//   assign u_8[183] = in_8[183] + e1_ext[2][183];
//   assign u_9[183] = in_9[183] + e1_ext[2][183];
//   assign u_1[184] = in_1[184] + e1_ext[0][184];
//   assign u_2[184] = in_2[184] + e1_ext[0][184];
//   assign u_3[184] = in_3[184] + e1_ext[0][184];
//   assign u_4[184] = in_4[184] + e1_ext[1][184];
//   assign u_5[184] = in_5[184] + e1_ext[1][184];
//   assign u_6[184] = in_6[184] + e1_ext[1][184];
//   assign u_7[184] = in_7[184] + e1_ext[2][184];
//   assign u_8[184] = in_8[184] + e1_ext[2][184];
//   assign u_9[184] = in_9[184] + e1_ext[2][184];
//   assign u_1[185] = in_1[185] + e1_ext[0][185];
//   assign u_2[185] = in_2[185] + e1_ext[0][185];
//   assign u_3[185] = in_3[185] + e1_ext[0][185];
//   assign u_4[185] = in_4[185] + e1_ext[1][185];
//   assign u_5[185] = in_5[185] + e1_ext[1][185];
//   assign u_6[185] = in_6[185] + e1_ext[1][185];
//   assign u_7[185] = in_7[185] + e1_ext[2][185];
//   assign u_8[185] = in_8[185] + e1_ext[2][185];
//   assign u_9[185] = in_9[185] + e1_ext[2][185];
//   assign u_1[186] = in_1[186] + e1_ext[0][186];
//   assign u_2[186] = in_2[186] + e1_ext[0][186];
//   assign u_3[186] = in_3[186] + e1_ext[0][186];
//   assign u_4[186] = in_4[186] + e1_ext[1][186];
//   assign u_5[186] = in_5[186] + e1_ext[1][186];
//   assign u_6[186] = in_6[186] + e1_ext[1][186];
//   assign u_7[186] = in_7[186] + e1_ext[2][186];
//   assign u_8[186] = in_8[186] + e1_ext[2][186];
//   assign u_9[186] = in_9[186] + e1_ext[2][186];
//   assign u_1[187] = in_1[187] + e1_ext[0][187];
//   assign u_2[187] = in_2[187] + e1_ext[0][187];
//   assign u_3[187] = in_3[187] + e1_ext[0][187];
//   assign u_4[187] = in_4[187] + e1_ext[1][187];
//   assign u_5[187] = in_5[187] + e1_ext[1][187];
//   assign u_6[187] = in_6[187] + e1_ext[1][187];
//   assign u_7[187] = in_7[187] + e1_ext[2][187];
//   assign u_8[187] = in_8[187] + e1_ext[2][187];
//   assign u_9[187] = in_9[187] + e1_ext[2][187];
//   assign u_1[188] = in_1[188] + e1_ext[0][188];
//   assign u_2[188] = in_2[188] + e1_ext[0][188];
//   assign u_3[188] = in_3[188] + e1_ext[0][188];
//   assign u_4[188] = in_4[188] + e1_ext[1][188];
//   assign u_5[188] = in_5[188] + e1_ext[1][188];
//   assign u_6[188] = in_6[188] + e1_ext[1][188];
//   assign u_7[188] = in_7[188] + e1_ext[2][188];
//   assign u_8[188] = in_8[188] + e1_ext[2][188];
//   assign u_9[188] = in_9[188] + e1_ext[2][188];
//   assign u_1[189] = in_1[189] + e1_ext[0][189];
//   assign u_2[189] = in_2[189] + e1_ext[0][189];
//   assign u_3[189] = in_3[189] + e1_ext[0][189];
//   assign u_4[189] = in_4[189] + e1_ext[1][189];
//   assign u_5[189] = in_5[189] + e1_ext[1][189];
//   assign u_6[189] = in_6[189] + e1_ext[1][189];
//   assign u_7[189] = in_7[189] + e1_ext[2][189];
//   assign u_8[189] = in_8[189] + e1_ext[2][189];
//   assign u_9[189] = in_9[189] + e1_ext[2][189];
//   assign u_1[190] = in_1[190] + e1_ext[0][190];
//   assign u_2[190] = in_2[190] + e1_ext[0][190];
//   assign u_3[190] = in_3[190] + e1_ext[0][190];
//   assign u_4[190] = in_4[190] + e1_ext[1][190];
//   assign u_5[190] = in_5[190] + e1_ext[1][190];
//   assign u_6[190] = in_6[190] + e1_ext[1][190];
//   assign u_7[190] = in_7[190] + e1_ext[2][190];
//   assign u_8[190] = in_8[190] + e1_ext[2][190];
//   assign u_9[190] = in_9[190] + e1_ext[2][190];
//   assign u_1[191] = in_1[191] + e1_ext[0][191];
//   assign u_2[191] = in_2[191] + e1_ext[0][191];
//   assign u_3[191] = in_3[191] + e1_ext[0][191];
//   assign u_4[191] = in_4[191] + e1_ext[1][191];
//   assign u_5[191] = in_5[191] + e1_ext[1][191];
//   assign u_6[191] = in_6[191] + e1_ext[1][191];
//   assign u_7[191] = in_7[191] + e1_ext[2][191];
//   assign u_8[191] = in_8[191] + e1_ext[2][191];
//   assign u_9[191] = in_9[191] + e1_ext[2][191];
//   assign u_1[192] = in_1[192] + e1_ext[0][192];
//   assign u_2[192] = in_2[192] + e1_ext[0][192];
//   assign u_3[192] = in_3[192] + e1_ext[0][192];
//   assign u_4[192] = in_4[192] + e1_ext[1][192];
//   assign u_5[192] = in_5[192] + e1_ext[1][192];
//   assign u_6[192] = in_6[192] + e1_ext[1][192];
//   assign u_7[192] = in_7[192] + e1_ext[2][192];
//   assign u_8[192] = in_8[192] + e1_ext[2][192];
//   assign u_9[192] = in_9[192] + e1_ext[2][192];
//   assign u_1[193] = in_1[193] + e1_ext[0][193];
//   assign u_2[193] = in_2[193] + e1_ext[0][193];
//   assign u_3[193] = in_3[193] + e1_ext[0][193];
//   assign u_4[193] = in_4[193] + e1_ext[1][193];
//   assign u_5[193] = in_5[193] + e1_ext[1][193];
//   assign u_6[193] = in_6[193] + e1_ext[1][193];
//   assign u_7[193] = in_7[193] + e1_ext[2][193];
//   assign u_8[193] = in_8[193] + e1_ext[2][193];
//   assign u_9[193] = in_9[193] + e1_ext[2][193];
//   assign u_1[194] = in_1[194] + e1_ext[0][194];
//   assign u_2[194] = in_2[194] + e1_ext[0][194];
//   assign u_3[194] = in_3[194] + e1_ext[0][194];
//   assign u_4[194] = in_4[194] + e1_ext[1][194];
//   assign u_5[194] = in_5[194] + e1_ext[1][194];
//   assign u_6[194] = in_6[194] + e1_ext[1][194];
//   assign u_7[194] = in_7[194] + e1_ext[2][194];
//   assign u_8[194] = in_8[194] + e1_ext[2][194];
//   assign u_9[194] = in_9[194] + e1_ext[2][194];
//   assign u_1[195] = in_1[195] + e1_ext[0][195];
//   assign u_2[195] = in_2[195] + e1_ext[0][195];
//   assign u_3[195] = in_3[195] + e1_ext[0][195];
//   assign u_4[195] = in_4[195] + e1_ext[1][195];
//   assign u_5[195] = in_5[195] + e1_ext[1][195];
//   assign u_6[195] = in_6[195] + e1_ext[1][195];
//   assign u_7[195] = in_7[195] + e1_ext[2][195];
//   assign u_8[195] = in_8[195] + e1_ext[2][195];
//   assign u_9[195] = in_9[195] + e1_ext[2][195];
//   assign u_1[196] = in_1[196] + e1_ext[0][196];
//   assign u_2[196] = in_2[196] + e1_ext[0][196];
//   assign u_3[196] = in_3[196] + e1_ext[0][196];
//   assign u_4[196] = in_4[196] + e1_ext[1][196];
//   assign u_5[196] = in_5[196] + e1_ext[1][196];
//   assign u_6[196] = in_6[196] + e1_ext[1][196];
//   assign u_7[196] = in_7[196] + e1_ext[2][196];
//   assign u_8[196] = in_8[196] + e1_ext[2][196];
//   assign u_9[196] = in_9[196] + e1_ext[2][196];
//   assign u_1[197] = in_1[197] + e1_ext[0][197];
//   assign u_2[197] = in_2[197] + e1_ext[0][197];
//   assign u_3[197] = in_3[197] + e1_ext[0][197];
//   assign u_4[197] = in_4[197] + e1_ext[1][197];
//   assign u_5[197] = in_5[197] + e1_ext[1][197];
//   assign u_6[197] = in_6[197] + e1_ext[1][197];
//   assign u_7[197] = in_7[197] + e1_ext[2][197];
//   assign u_8[197] = in_8[197] + e1_ext[2][197];
//   assign u_9[197] = in_9[197] + e1_ext[2][197];
//   assign u_1[198] = in_1[198] + e1_ext[0][198];
//   assign u_2[198] = in_2[198] + e1_ext[0][198];
//   assign u_3[198] = in_3[198] + e1_ext[0][198];
//   assign u_4[198] = in_4[198] + e1_ext[1][198];
//   assign u_5[198] = in_5[198] + e1_ext[1][198];
//   assign u_6[198] = in_6[198] + e1_ext[1][198];
//   assign u_7[198] = in_7[198] + e1_ext[2][198];
//   assign u_8[198] = in_8[198] + e1_ext[2][198];
//   assign u_9[198] = in_9[198] + e1_ext[2][198];
//   assign u_1[199] = in_1[199] + e1_ext[0][199];
//   assign u_2[199] = in_2[199] + e1_ext[0][199];
//   assign u_3[199] = in_3[199] + e1_ext[0][199];
//   assign u_4[199] = in_4[199] + e1_ext[1][199];
//   assign u_5[199] = in_5[199] + e1_ext[1][199];
//   assign u_6[199] = in_6[199] + e1_ext[1][199];
//   assign u_7[199] = in_7[199] + e1_ext[2][199];
//   assign u_8[199] = in_8[199] + e1_ext[2][199];
//   assign u_9[199] = in_9[199] + e1_ext[2][199];
//   assign u_1[200] = in_1[200] + e1_ext[0][200];
//   assign u_2[200] = in_2[200] + e1_ext[0][200];
//   assign u_3[200] = in_3[200] + e1_ext[0][200];
//   assign u_4[200] = in_4[200] + e1_ext[1][200];
//   assign u_5[200] = in_5[200] + e1_ext[1][200];
//   assign u_6[200] = in_6[200] + e1_ext[1][200];
//   assign u_7[200] = in_7[200] + e1_ext[2][200];
//   assign u_8[200] = in_8[200] + e1_ext[2][200];
//   assign u_9[200] = in_9[200] + e1_ext[2][200];
//   assign u_1[201] = in_1[201] + e1_ext[0][201];
//   assign u_2[201] = in_2[201] + e1_ext[0][201];
//   assign u_3[201] = in_3[201] + e1_ext[0][201];
//   assign u_4[201] = in_4[201] + e1_ext[1][201];
//   assign u_5[201] = in_5[201] + e1_ext[1][201];
//   assign u_6[201] = in_6[201] + e1_ext[1][201];
//   assign u_7[201] = in_7[201] + e1_ext[2][201];
//   assign u_8[201] = in_8[201] + e1_ext[2][201];
//   assign u_9[201] = in_9[201] + e1_ext[2][201];
//   assign u_1[202] = in_1[202] + e1_ext[0][202];
//   assign u_2[202] = in_2[202] + e1_ext[0][202];
//   assign u_3[202] = in_3[202] + e1_ext[0][202];
//   assign u_4[202] = in_4[202] + e1_ext[1][202];
//   assign u_5[202] = in_5[202] + e1_ext[1][202];
//   assign u_6[202] = in_6[202] + e1_ext[1][202];
//   assign u_7[202] = in_7[202] + e1_ext[2][202];
//   assign u_8[202] = in_8[202] + e1_ext[2][202];
//   assign u_9[202] = in_9[202] + e1_ext[2][202];
//   assign u_1[203] = in_1[203] + e1_ext[0][203];
//   assign u_2[203] = in_2[203] + e1_ext[0][203];
//   assign u_3[203] = in_3[203] + e1_ext[0][203];
//   assign u_4[203] = in_4[203] + e1_ext[1][203];
//   assign u_5[203] = in_5[203] + e1_ext[1][203];
//   assign u_6[203] = in_6[203] + e1_ext[1][203];
//   assign u_7[203] = in_7[203] + e1_ext[2][203];
//   assign u_8[203] = in_8[203] + e1_ext[2][203];
//   assign u_9[203] = in_9[203] + e1_ext[2][203];
//   assign u_1[204] = in_1[204] + e1_ext[0][204];
//   assign u_2[204] = in_2[204] + e1_ext[0][204];
//   assign u_3[204] = in_3[204] + e1_ext[0][204];
//   assign u_4[204] = in_4[204] + e1_ext[1][204];
//   assign u_5[204] = in_5[204] + e1_ext[1][204];
//   assign u_6[204] = in_6[204] + e1_ext[1][204];
//   assign u_7[204] = in_7[204] + e1_ext[2][204];
//   assign u_8[204] = in_8[204] + e1_ext[2][204];
//   assign u_9[204] = in_9[204] + e1_ext[2][204];
//   assign u_1[205] = in_1[205] + e1_ext[0][205];
//   assign u_2[205] = in_2[205] + e1_ext[0][205];
//   assign u_3[205] = in_3[205] + e1_ext[0][205];
//   assign u_4[205] = in_4[205] + e1_ext[1][205];
//   assign u_5[205] = in_5[205] + e1_ext[1][205];
//   assign u_6[205] = in_6[205] + e1_ext[1][205];
//   assign u_7[205] = in_7[205] + e1_ext[2][205];
//   assign u_8[205] = in_8[205] + e1_ext[2][205];
//   assign u_9[205] = in_9[205] + e1_ext[2][205];
//   assign u_1[206] = in_1[206] + e1_ext[0][206];
//   assign u_2[206] = in_2[206] + e1_ext[0][206];
//   assign u_3[206] = in_3[206] + e1_ext[0][206];
//   assign u_4[206] = in_4[206] + e1_ext[1][206];
//   assign u_5[206] = in_5[206] + e1_ext[1][206];
//   assign u_6[206] = in_6[206] + e1_ext[1][206];
//   assign u_7[206] = in_7[206] + e1_ext[2][206];
//   assign u_8[206] = in_8[206] + e1_ext[2][206];
//   assign u_9[206] = in_9[206] + e1_ext[2][206];
//   assign u_1[207] = in_1[207] + e1_ext[0][207];
//   assign u_2[207] = in_2[207] + e1_ext[0][207];
//   assign u_3[207] = in_3[207] + e1_ext[0][207];
//   assign u_4[207] = in_4[207] + e1_ext[1][207];
//   assign u_5[207] = in_5[207] + e1_ext[1][207];
//   assign u_6[207] = in_6[207] + e1_ext[1][207];
//   assign u_7[207] = in_7[207] + e1_ext[2][207];
//   assign u_8[207] = in_8[207] + e1_ext[2][207];
//   assign u_9[207] = in_9[207] + e1_ext[2][207];
//   assign u_1[208] = in_1[208] + e1_ext[0][208];
//   assign u_2[208] = in_2[208] + e1_ext[0][208];
//   assign u_3[208] = in_3[208] + e1_ext[0][208];
//   assign u_4[208] = in_4[208] + e1_ext[1][208];
//   assign u_5[208] = in_5[208] + e1_ext[1][208];
//   assign u_6[208] = in_6[208] + e1_ext[1][208];
//   assign u_7[208] = in_7[208] + e1_ext[2][208];
//   assign u_8[208] = in_8[208] + e1_ext[2][208];
//   assign u_9[208] = in_9[208] + e1_ext[2][208];
//   assign u_1[209] = in_1[209] + e1_ext[0][209];
//   assign u_2[209] = in_2[209] + e1_ext[0][209];
//   assign u_3[209] = in_3[209] + e1_ext[0][209];
//   assign u_4[209] = in_4[209] + e1_ext[1][209];
//   assign u_5[209] = in_5[209] + e1_ext[1][209];
//   assign u_6[209] = in_6[209] + e1_ext[1][209];
//   assign u_7[209] = in_7[209] + e1_ext[2][209];
//   assign u_8[209] = in_8[209] + e1_ext[2][209];
//   assign u_9[209] = in_9[209] + e1_ext[2][209];
//   assign u_1[210] = in_1[210] + e1_ext[0][210];
//   assign u_2[210] = in_2[210] + e1_ext[0][210];
//   assign u_3[210] = in_3[210] + e1_ext[0][210];
//   assign u_4[210] = in_4[210] + e1_ext[1][210];
//   assign u_5[210] = in_5[210] + e1_ext[1][210];
//   assign u_6[210] = in_6[210] + e1_ext[1][210];
//   assign u_7[210] = in_7[210] + e1_ext[2][210];
//   assign u_8[210] = in_8[210] + e1_ext[2][210];
//   assign u_9[210] = in_9[210] + e1_ext[2][210];
//   assign u_1[211] = in_1[211] + e1_ext[0][211];
//   assign u_2[211] = in_2[211] + e1_ext[0][211];
//   assign u_3[211] = in_3[211] + e1_ext[0][211];
//   assign u_4[211] = in_4[211] + e1_ext[1][211];
//   assign u_5[211] = in_5[211] + e1_ext[1][211];
//   assign u_6[211] = in_6[211] + e1_ext[1][211];
//   assign u_7[211] = in_7[211] + e1_ext[2][211];
//   assign u_8[211] = in_8[211] + e1_ext[2][211];
//   assign u_9[211] = in_9[211] + e1_ext[2][211];
//   assign u_1[212] = in_1[212] + e1_ext[0][212];
//   assign u_2[212] = in_2[212] + e1_ext[0][212];
//   assign u_3[212] = in_3[212] + e1_ext[0][212];
//   assign u_4[212] = in_4[212] + e1_ext[1][212];
//   assign u_5[212] = in_5[212] + e1_ext[1][212];
//   assign u_6[212] = in_6[212] + e1_ext[1][212];
//   assign u_7[212] = in_7[212] + e1_ext[2][212];
//   assign u_8[212] = in_8[212] + e1_ext[2][212];
//   assign u_9[212] = in_9[212] + e1_ext[2][212];
//   assign u_1[213] = in_1[213] + e1_ext[0][213];
//   assign u_2[213] = in_2[213] + e1_ext[0][213];
//   assign u_3[213] = in_3[213] + e1_ext[0][213];
//   assign u_4[213] = in_4[213] + e1_ext[1][213];
//   assign u_5[213] = in_5[213] + e1_ext[1][213];
//   assign u_6[213] = in_6[213] + e1_ext[1][213];
//   assign u_7[213] = in_7[213] + e1_ext[2][213];
//   assign u_8[213] = in_8[213] + e1_ext[2][213];
//   assign u_9[213] = in_9[213] + e1_ext[2][213];
//   assign u_1[214] = in_1[214] + e1_ext[0][214];
//   assign u_2[214] = in_2[214] + e1_ext[0][214];
//   assign u_3[214] = in_3[214] + e1_ext[0][214];
//   assign u_4[214] = in_4[214] + e1_ext[1][214];
//   assign u_5[214] = in_5[214] + e1_ext[1][214];
//   assign u_6[214] = in_6[214] + e1_ext[1][214];
//   assign u_7[214] = in_7[214] + e1_ext[2][214];
//   assign u_8[214] = in_8[214] + e1_ext[2][214];
//   assign u_9[214] = in_9[214] + e1_ext[2][214];
//   assign u_1[215] = in_1[215] + e1_ext[0][215];
//   assign u_2[215] = in_2[215] + e1_ext[0][215];
//   assign u_3[215] = in_3[215] + e1_ext[0][215];
//   assign u_4[215] = in_4[215] + e1_ext[1][215];
//   assign u_5[215] = in_5[215] + e1_ext[1][215];
//   assign u_6[215] = in_6[215] + e1_ext[1][215];
//   assign u_7[215] = in_7[215] + e1_ext[2][215];
//   assign u_8[215] = in_8[215] + e1_ext[2][215];
//   assign u_9[215] = in_9[215] + e1_ext[2][215];
//   assign u_1[216] = in_1[216] + e1_ext[0][216];
//   assign u_2[216] = in_2[216] + e1_ext[0][216];
//   assign u_3[216] = in_3[216] + e1_ext[0][216];
//   assign u_4[216] = in_4[216] + e1_ext[1][216];
//   assign u_5[216] = in_5[216] + e1_ext[1][216];
//   assign u_6[216] = in_6[216] + e1_ext[1][216];
//   assign u_7[216] = in_7[216] + e1_ext[2][216];
//   assign u_8[216] = in_8[216] + e1_ext[2][216];
//   assign u_9[216] = in_9[216] + e1_ext[2][216];
//   assign u_1[217] = in_1[217] + e1_ext[0][217];
//   assign u_2[217] = in_2[217] + e1_ext[0][217];
//   assign u_3[217] = in_3[217] + e1_ext[0][217];
//   assign u_4[217] = in_4[217] + e1_ext[1][217];
//   assign u_5[217] = in_5[217] + e1_ext[1][217];
//   assign u_6[217] = in_6[217] + e1_ext[1][217];
//   assign u_7[217] = in_7[217] + e1_ext[2][217];
//   assign u_8[217] = in_8[217] + e1_ext[2][217];
//   assign u_9[217] = in_9[217] + e1_ext[2][217];
//   assign u_1[218] = in_1[218] + e1_ext[0][218];
//   assign u_2[218] = in_2[218] + e1_ext[0][218];
//   assign u_3[218] = in_3[218] + e1_ext[0][218];
//   assign u_4[218] = in_4[218] + e1_ext[1][218];
//   assign u_5[218] = in_5[218] + e1_ext[1][218];
//   assign u_6[218] = in_6[218] + e1_ext[1][218];
//   assign u_7[218] = in_7[218] + e1_ext[2][218];
//   assign u_8[218] = in_8[218] + e1_ext[2][218];
//   assign u_9[218] = in_9[218] + e1_ext[2][218];
//   assign u_1[219] = in_1[219] + e1_ext[0][219];
//   assign u_2[219] = in_2[219] + e1_ext[0][219];
//   assign u_3[219] = in_3[219] + e1_ext[0][219];
//   assign u_4[219] = in_4[219] + e1_ext[1][219];
//   assign u_5[219] = in_5[219] + e1_ext[1][219];
//   assign u_6[219] = in_6[219] + e1_ext[1][219];
//   assign u_7[219] = in_7[219] + e1_ext[2][219];
//   assign u_8[219] = in_8[219] + e1_ext[2][219];
//   assign u_9[219] = in_9[219] + e1_ext[2][219];
//   assign u_1[220] = in_1[220] + e1_ext[0][220];
//   assign u_2[220] = in_2[220] + e1_ext[0][220];
//   assign u_3[220] = in_3[220] + e1_ext[0][220];
//   assign u_4[220] = in_4[220] + e1_ext[1][220];
//   assign u_5[220] = in_5[220] + e1_ext[1][220];
//   assign u_6[220] = in_6[220] + e1_ext[1][220];
//   assign u_7[220] = in_7[220] + e1_ext[2][220];
//   assign u_8[220] = in_8[220] + e1_ext[2][220];
//   assign u_9[220] = in_9[220] + e1_ext[2][220];
//   assign u_1[221] = in_1[221] + e1_ext[0][221];
//   assign u_2[221] = in_2[221] + e1_ext[0][221];
//   assign u_3[221] = in_3[221] + e1_ext[0][221];
//   assign u_4[221] = in_4[221] + e1_ext[1][221];
//   assign u_5[221] = in_5[221] + e1_ext[1][221];
//   assign u_6[221] = in_6[221] + e1_ext[1][221];
//   assign u_7[221] = in_7[221] + e1_ext[2][221];
//   assign u_8[221] = in_8[221] + e1_ext[2][221];
//   assign u_9[221] = in_9[221] + e1_ext[2][221];
//   assign u_1[222] = in_1[222] + e1_ext[0][222];
//   assign u_2[222] = in_2[222] + e1_ext[0][222];
//   assign u_3[222] = in_3[222] + e1_ext[0][222];
//   assign u_4[222] = in_4[222] + e1_ext[1][222];
//   assign u_5[222] = in_5[222] + e1_ext[1][222];
//   assign u_6[222] = in_6[222] + e1_ext[1][222];
//   assign u_7[222] = in_7[222] + e1_ext[2][222];
//   assign u_8[222] = in_8[222] + e1_ext[2][222];
//   assign u_9[222] = in_9[222] + e1_ext[2][222];
//   assign u_1[223] = in_1[223] + e1_ext[0][223];
//   assign u_2[223] = in_2[223] + e1_ext[0][223];
//   assign u_3[223] = in_3[223] + e1_ext[0][223];
//   assign u_4[223] = in_4[223] + e1_ext[1][223];
//   assign u_5[223] = in_5[223] + e1_ext[1][223];
//   assign u_6[223] = in_6[223] + e1_ext[1][223];
//   assign u_7[223] = in_7[223] + e1_ext[2][223];
//   assign u_8[223] = in_8[223] + e1_ext[2][223];
//   assign u_9[223] = in_9[223] + e1_ext[2][223];
//   assign u_1[224] = in_1[224] + e1_ext[0][224];
//   assign u_2[224] = in_2[224] + e1_ext[0][224];
//   assign u_3[224] = in_3[224] + e1_ext[0][224];
//   assign u_4[224] = in_4[224] + e1_ext[1][224];
//   assign u_5[224] = in_5[224] + e1_ext[1][224];
//   assign u_6[224] = in_6[224] + e1_ext[1][224];
//   assign u_7[224] = in_7[224] + e1_ext[2][224];
//   assign u_8[224] = in_8[224] + e1_ext[2][224];
//   assign u_9[224] = in_9[224] + e1_ext[2][224];
//   assign u_1[225] = in_1[225] + e1_ext[0][225];
//   assign u_2[225] = in_2[225] + e1_ext[0][225];
//   assign u_3[225] = in_3[225] + e1_ext[0][225];
//   assign u_4[225] = in_4[225] + e1_ext[1][225];
//   assign u_5[225] = in_5[225] + e1_ext[1][225];
//   assign u_6[225] = in_6[225] + e1_ext[1][225];
//   assign u_7[225] = in_7[225] + e1_ext[2][225];
//   assign u_8[225] = in_8[225] + e1_ext[2][225];
//   assign u_9[225] = in_9[225] + e1_ext[2][225];
//   assign u_1[226] = in_1[226] + e1_ext[0][226];
//   assign u_2[226] = in_2[226] + e1_ext[0][226];
//   assign u_3[226] = in_3[226] + e1_ext[0][226];
//   assign u_4[226] = in_4[226] + e1_ext[1][226];
//   assign u_5[226] = in_5[226] + e1_ext[1][226];
//   assign u_6[226] = in_6[226] + e1_ext[1][226];
//   assign u_7[226] = in_7[226] + e1_ext[2][226];
//   assign u_8[226] = in_8[226] + e1_ext[2][226];
//   assign u_9[226] = in_9[226] + e1_ext[2][226];
//   assign u_1[227] = in_1[227] + e1_ext[0][227];
//   assign u_2[227] = in_2[227] + e1_ext[0][227];
//   assign u_3[227] = in_3[227] + e1_ext[0][227];
//   assign u_4[227] = in_4[227] + e1_ext[1][227];
//   assign u_5[227] = in_5[227] + e1_ext[1][227];
//   assign u_6[227] = in_6[227] + e1_ext[1][227];
//   assign u_7[227] = in_7[227] + e1_ext[2][227];
//   assign u_8[227] = in_8[227] + e1_ext[2][227];
//   assign u_9[227] = in_9[227] + e1_ext[2][227];
//   assign u_1[228] = in_1[228] + e1_ext[0][228];
//   assign u_2[228] = in_2[228] + e1_ext[0][228];
//   assign u_3[228] = in_3[228] + e1_ext[0][228];
//   assign u_4[228] = in_4[228] + e1_ext[1][228];
//   assign u_5[228] = in_5[228] + e1_ext[1][228];
//   assign u_6[228] = in_6[228] + e1_ext[1][228];
//   assign u_7[228] = in_7[228] + e1_ext[2][228];
//   assign u_8[228] = in_8[228] + e1_ext[2][228];
//   assign u_9[228] = in_9[228] + e1_ext[2][228];
//   assign u_1[229] = in_1[229] + e1_ext[0][229];
//   assign u_2[229] = in_2[229] + e1_ext[0][229];
//   assign u_3[229] = in_3[229] + e1_ext[0][229];
//   assign u_4[229] = in_4[229] + e1_ext[1][229];
//   assign u_5[229] = in_5[229] + e1_ext[1][229];
//   assign u_6[229] = in_6[229] + e1_ext[1][229];
//   assign u_7[229] = in_7[229] + e1_ext[2][229];
//   assign u_8[229] = in_8[229] + e1_ext[2][229];
//   assign u_9[229] = in_9[229] + e1_ext[2][229];
//   assign u_1[230] = in_1[230] + e1_ext[0][230];
//   assign u_2[230] = in_2[230] + e1_ext[0][230];
//   assign u_3[230] = in_3[230] + e1_ext[0][230];
//   assign u_4[230] = in_4[230] + e1_ext[1][230];
//   assign u_5[230] = in_5[230] + e1_ext[1][230];
//   assign u_6[230] = in_6[230] + e1_ext[1][230];
//   assign u_7[230] = in_7[230] + e1_ext[2][230];
//   assign u_8[230] = in_8[230] + e1_ext[2][230];
//   assign u_9[230] = in_9[230] + e1_ext[2][230];
//   assign u_1[231] = in_1[231] + e1_ext[0][231];
//   assign u_2[231] = in_2[231] + e1_ext[0][231];
//   assign u_3[231] = in_3[231] + e1_ext[0][231];
//   assign u_4[231] = in_4[231] + e1_ext[1][231];
//   assign u_5[231] = in_5[231] + e1_ext[1][231];
//   assign u_6[231] = in_6[231] + e1_ext[1][231];
//   assign u_7[231] = in_7[231] + e1_ext[2][231];
//   assign u_8[231] = in_8[231] + e1_ext[2][231];
//   assign u_9[231] = in_9[231] + e1_ext[2][231];
//   assign u_1[232] = in_1[232] + e1_ext[0][232];
//   assign u_2[232] = in_2[232] + e1_ext[0][232];
//   assign u_3[232] = in_3[232] + e1_ext[0][232];
//   assign u_4[232] = in_4[232] + e1_ext[1][232];
//   assign u_5[232] = in_5[232] + e1_ext[1][232];
//   assign u_6[232] = in_6[232] + e1_ext[1][232];
//   assign u_7[232] = in_7[232] + e1_ext[2][232];
//   assign u_8[232] = in_8[232] + e1_ext[2][232];
//   assign u_9[232] = in_9[232] + e1_ext[2][232];
//   assign u_1[233] = in_1[233] + e1_ext[0][233];
//   assign u_2[233] = in_2[233] + e1_ext[0][233];
//   assign u_3[233] = in_3[233] + e1_ext[0][233];
//   assign u_4[233] = in_4[233] + e1_ext[1][233];
//   assign u_5[233] = in_5[233] + e1_ext[1][233];
//   assign u_6[233] = in_6[233] + e1_ext[1][233];
//   assign u_7[233] = in_7[233] + e1_ext[2][233];
//   assign u_8[233] = in_8[233] + e1_ext[2][233];
//   assign u_9[233] = in_9[233] + e1_ext[2][233];
//   assign u_1[234] = in_1[234] + e1_ext[0][234];
//   assign u_2[234] = in_2[234] + e1_ext[0][234];
//   assign u_3[234] = in_3[234] + e1_ext[0][234];
//   assign u_4[234] = in_4[234] + e1_ext[1][234];
//   assign u_5[234] = in_5[234] + e1_ext[1][234];
//   assign u_6[234] = in_6[234] + e1_ext[1][234];
//   assign u_7[234] = in_7[234] + e1_ext[2][234];
//   assign u_8[234] = in_8[234] + e1_ext[2][234];
//   assign u_9[234] = in_9[234] + e1_ext[2][234];
//   assign u_1[235] = in_1[235] + e1_ext[0][235];
//   assign u_2[235] = in_2[235] + e1_ext[0][235];
//   assign u_3[235] = in_3[235] + e1_ext[0][235];
//   assign u_4[235] = in_4[235] + e1_ext[1][235];
//   assign u_5[235] = in_5[235] + e1_ext[1][235];
//   assign u_6[235] = in_6[235] + e1_ext[1][235];
//   assign u_7[235] = in_7[235] + e1_ext[2][235];
//   assign u_8[235] = in_8[235] + e1_ext[2][235];
//   assign u_9[235] = in_9[235] + e1_ext[2][235];
//   assign u_1[236] = in_1[236] + e1_ext[0][236];
//   assign u_2[236] = in_2[236] + e1_ext[0][236];
//   assign u_3[236] = in_3[236] + e1_ext[0][236];
//   assign u_4[236] = in_4[236] + e1_ext[1][236];
//   assign u_5[236] = in_5[236] + e1_ext[1][236];
//   assign u_6[236] = in_6[236] + e1_ext[1][236];
//   assign u_7[236] = in_7[236] + e1_ext[2][236];
//   assign u_8[236] = in_8[236] + e1_ext[2][236];
//   assign u_9[236] = in_9[236] + e1_ext[2][236];
//   assign u_1[237] = in_1[237] + e1_ext[0][237];
//   assign u_2[237] = in_2[237] + e1_ext[0][237];
//   assign u_3[237] = in_3[237] + e1_ext[0][237];
//   assign u_4[237] = in_4[237] + e1_ext[1][237];
//   assign u_5[237] = in_5[237] + e1_ext[1][237];
//   assign u_6[237] = in_6[237] + e1_ext[1][237];
//   assign u_7[237] = in_7[237] + e1_ext[2][237];
//   assign u_8[237] = in_8[237] + e1_ext[2][237];
//   assign u_9[237] = in_9[237] + e1_ext[2][237];
//   assign u_1[238] = in_1[238] + e1_ext[0][238];
//   assign u_2[238] = in_2[238] + e1_ext[0][238];
//   assign u_3[238] = in_3[238] + e1_ext[0][238];
//   assign u_4[238] = in_4[238] + e1_ext[1][238];
//   assign u_5[238] = in_5[238] + e1_ext[1][238];
//   assign u_6[238] = in_6[238] + e1_ext[1][238];
//   assign u_7[238] = in_7[238] + e1_ext[2][238];
//   assign u_8[238] = in_8[238] + e1_ext[2][238];
//   assign u_9[238] = in_9[238] + e1_ext[2][238];
//   assign u_1[239] = in_1[239] + e1_ext[0][239];
//   assign u_2[239] = in_2[239] + e1_ext[0][239];
//   assign u_3[239] = in_3[239] + e1_ext[0][239];
//   assign u_4[239] = in_4[239] + e1_ext[1][239];
//   assign u_5[239] = in_5[239] + e1_ext[1][239];
//   assign u_6[239] = in_6[239] + e1_ext[1][239];
//   assign u_7[239] = in_7[239] + e1_ext[2][239];
//   assign u_8[239] = in_8[239] + e1_ext[2][239];
//   assign u_9[239] = in_9[239] + e1_ext[2][239];
//   assign u_1[240] = in_1[240] + e1_ext[0][240];
//   assign u_2[240] = in_2[240] + e1_ext[0][240];
//   assign u_3[240] = in_3[240] + e1_ext[0][240];
//   assign u_4[240] = in_4[240] + e1_ext[1][240];
//   assign u_5[240] = in_5[240] + e1_ext[1][240];
//   assign u_6[240] = in_6[240] + e1_ext[1][240];
//   assign u_7[240] = in_7[240] + e1_ext[2][240];
//   assign u_8[240] = in_8[240] + e1_ext[2][240];
//   assign u_9[240] = in_9[240] + e1_ext[2][240];
//   assign u_1[241] = in_1[241] + e1_ext[0][241];
//   assign u_2[241] = in_2[241] + e1_ext[0][241];
//   assign u_3[241] = in_3[241] + e1_ext[0][241];
//   assign u_4[241] = in_4[241] + e1_ext[1][241];
//   assign u_5[241] = in_5[241] + e1_ext[1][241];
//   assign u_6[241] = in_6[241] + e1_ext[1][241];
//   assign u_7[241] = in_7[241] + e1_ext[2][241];
//   assign u_8[241] = in_8[241] + e1_ext[2][241];
//   assign u_9[241] = in_9[241] + e1_ext[2][241];
//   assign u_1[242] = in_1[242] + e1_ext[0][242];
//   assign u_2[242] = in_2[242] + e1_ext[0][242];
//   assign u_3[242] = in_3[242] + e1_ext[0][242];
//   assign u_4[242] = in_4[242] + e1_ext[1][242];
//   assign u_5[242] = in_5[242] + e1_ext[1][242];
//   assign u_6[242] = in_6[242] + e1_ext[1][242];
//   assign u_7[242] = in_7[242] + e1_ext[2][242];
//   assign u_8[242] = in_8[242] + e1_ext[2][242];
//   assign u_9[242] = in_9[242] + e1_ext[2][242];
//   assign u_1[243] = in_1[243] + e1_ext[0][243];
//   assign u_2[243] = in_2[243] + e1_ext[0][243];
//   assign u_3[243] = in_3[243] + e1_ext[0][243];
//   assign u_4[243] = in_4[243] + e1_ext[1][243];
//   assign u_5[243] = in_5[243] + e1_ext[1][243];
//   assign u_6[243] = in_6[243] + e1_ext[1][243];
//   assign u_7[243] = in_7[243] + e1_ext[2][243];
//   assign u_8[243] = in_8[243] + e1_ext[2][243];
//   assign u_9[243] = in_9[243] + e1_ext[2][243];
//   assign u_1[244] = in_1[244] + e1_ext[0][244];
//   assign u_2[244] = in_2[244] + e1_ext[0][244];
//   assign u_3[244] = in_3[244] + e1_ext[0][244];
//   assign u_4[244] = in_4[244] + e1_ext[1][244];
//   assign u_5[244] = in_5[244] + e1_ext[1][244];
//   assign u_6[244] = in_6[244] + e1_ext[1][244];
//   assign u_7[244] = in_7[244] + e1_ext[2][244];
//   assign u_8[244] = in_8[244] + e1_ext[2][244];
//   assign u_9[244] = in_9[244] + e1_ext[2][244];
//   assign u_1[245] = in_1[245] + e1_ext[0][245];
//   assign u_2[245] = in_2[245] + e1_ext[0][245];
//   assign u_3[245] = in_3[245] + e1_ext[0][245];
//   assign u_4[245] = in_4[245] + e1_ext[1][245];
//   assign u_5[245] = in_5[245] + e1_ext[1][245];
//   assign u_6[245] = in_6[245] + e1_ext[1][245];
//   assign u_7[245] = in_7[245] + e1_ext[2][245];
//   assign u_8[245] = in_8[245] + e1_ext[2][245];
//   assign u_9[245] = in_9[245] + e1_ext[2][245];
//   assign u_1[246] = in_1[246] + e1_ext[0][246];
//   assign u_2[246] = in_2[246] + e1_ext[0][246];
//   assign u_3[246] = in_3[246] + e1_ext[0][246];
//   assign u_4[246] = in_4[246] + e1_ext[1][246];
//   assign u_5[246] = in_5[246] + e1_ext[1][246];
//   assign u_6[246] = in_6[246] + e1_ext[1][246];
//   assign u_7[246] = in_7[246] + e1_ext[2][246];
//   assign u_8[246] = in_8[246] + e1_ext[2][246];
//   assign u_9[246] = in_9[246] + e1_ext[2][246];
//   assign u_1[247] = in_1[247] + e1_ext[0][247];
//   assign u_2[247] = in_2[247] + e1_ext[0][247];
//   assign u_3[247] = in_3[247] + e1_ext[0][247];
//   assign u_4[247] = in_4[247] + e1_ext[1][247];
//   assign u_5[247] = in_5[247] + e1_ext[1][247];
//   assign u_6[247] = in_6[247] + e1_ext[1][247];
//   assign u_7[247] = in_7[247] + e1_ext[2][247];
//   assign u_8[247] = in_8[247] + e1_ext[2][247];
//   assign u_9[247] = in_9[247] + e1_ext[2][247];
//   assign u_1[248] = in_1[248] + e1_ext[0][248];
//   assign u_2[248] = in_2[248] + e1_ext[0][248];
//   assign u_3[248] = in_3[248] + e1_ext[0][248];
//   assign u_4[248] = in_4[248] + e1_ext[1][248];
//   assign u_5[248] = in_5[248] + e1_ext[1][248];
//   assign u_6[248] = in_6[248] + e1_ext[1][248];
//   assign u_7[248] = in_7[248] + e1_ext[2][248];
//   assign u_8[248] = in_8[248] + e1_ext[2][248];
//   assign u_9[248] = in_9[248] + e1_ext[2][248];
//   assign u_1[249] = in_1[249] + e1_ext[0][249];
//   assign u_2[249] = in_2[249] + e1_ext[0][249];
//   assign u_3[249] = in_3[249] + e1_ext[0][249];
//   assign u_4[249] = in_4[249] + e1_ext[1][249];
//   assign u_5[249] = in_5[249] + e1_ext[1][249];
//   assign u_6[249] = in_6[249] + e1_ext[1][249];
//   assign u_7[249] = in_7[249] + e1_ext[2][249];
//   assign u_8[249] = in_8[249] + e1_ext[2][249];
//   assign u_9[249] = in_9[249] + e1_ext[2][249];
//   assign u_1[250] = in_1[250] + e1_ext[0][250];
//   assign u_2[250] = in_2[250] + e1_ext[0][250];
//   assign u_3[250] = in_3[250] + e1_ext[0][250];
//   assign u_4[250] = in_4[250] + e1_ext[1][250];
//   assign u_5[250] = in_5[250] + e1_ext[1][250];
//   assign u_6[250] = in_6[250] + e1_ext[1][250];
//   assign u_7[250] = in_7[250] + e1_ext[2][250];
//   assign u_8[250] = in_8[250] + e1_ext[2][250];
//   assign u_9[250] = in_9[250] + e1_ext[2][250];
//   assign u_1[251] = in_1[251] + e1_ext[0][251];
//   assign u_2[251] = in_2[251] + e1_ext[0][251];
//   assign u_3[251] = in_3[251] + e1_ext[0][251];
//   assign u_4[251] = in_4[251] + e1_ext[1][251];
//   assign u_5[251] = in_5[251] + e1_ext[1][251];
//   assign u_6[251] = in_6[251] + e1_ext[1][251];
//   assign u_7[251] = in_7[251] + e1_ext[2][251];
//   assign u_8[251] = in_8[251] + e1_ext[2][251];
//   assign u_9[251] = in_9[251] + e1_ext[2][251];
//   assign u_1[252] = in_1[252] + e1_ext[0][252];
//   assign u_2[252] = in_2[252] + e1_ext[0][252];
//   assign u_3[252] = in_3[252] + e1_ext[0][252];
//   assign u_4[252] = in_4[252] + e1_ext[1][252];
//   assign u_5[252] = in_5[252] + e1_ext[1][252];
//   assign u_6[252] = in_6[252] + e1_ext[1][252];
//   assign u_7[252] = in_7[252] + e1_ext[2][252];
//   assign u_8[252] = in_8[252] + e1_ext[2][252];
//   assign u_9[252] = in_9[252] + e1_ext[2][252];
//   assign u_1[253] = in_1[253] + e1_ext[0][253];
//   assign u_2[253] = in_2[253] + e1_ext[0][253];
//   assign u_3[253] = in_3[253] + e1_ext[0][253];
//   assign u_4[253] = in_4[253] + e1_ext[1][253];
//   assign u_5[253] = in_5[253] + e1_ext[1][253];
//   assign u_6[253] = in_6[253] + e1_ext[1][253];
//   assign u_7[253] = in_7[253] + e1_ext[2][253];
//   assign u_8[253] = in_8[253] + e1_ext[2][253];
//   assign u_9[253] = in_9[253] + e1_ext[2][253];
//   assign u_1[254] = in_1[254] + e1_ext[0][254];
//   assign u_2[254] = in_2[254] + e1_ext[0][254];
//   assign u_3[254] = in_3[254] + e1_ext[0][254];
//   assign u_4[254] = in_4[254] + e1_ext[1][254];
//   assign u_5[254] = in_5[254] + e1_ext[1][254];
//   assign u_6[254] = in_6[254] + e1_ext[1][254];
//   assign u_7[254] = in_7[254] + e1_ext[2][254];
//   assign u_8[254] = in_8[254] + e1_ext[2][254];
//   assign u_9[254] = in_9[254] + e1_ext[2][254];
//   assign u_1[255] = in_1[255] + e1_ext[0][255];
//   assign u_2[255] = in_2[255] + e1_ext[0][255];
//   assign u_3[255] = in_3[255] + e1_ext[0][255];
//   assign u_4[255] = in_4[255] + e1_ext[1][255];
//   assign u_5[255] = in_5[255] + e1_ext[1][255];
//   assign u_6[255] = in_6[255] + e1_ext[1][255];
//   assign u_7[255] = in_7[255] + e1_ext[2][255];
//   assign u_8[255] = in_8[255] + e1_ext[2][255];
//   assign u_9[255] = in_9[255] + e1_ext[2][255];



////assign m_slice0 = m[38:0];

// decode #(.ELL(16), .NUM_COEFFS(256), .BYTE_COUNT(32)) dec4 (
//       .byte_array(m),
//       .len(32),
//       .coeffs(m_dec)
//   );
   


//decompress_module decompress_inst0 (
//    .x(16),
//    .d(m_dec[0]),
//    .result(decom_out[0])
//);

//decompress_module decompress_inst1 (
//    .x(16),
//    .d(m_dec[1]),
//    .result(decom_out[1])
//);

//decompress_module decompress_inst2 (
//    .x(16),
//    .d(m_dec[2]),
//    .result(decom_out[2])
//);

//decompress_module decompress_inst3 (
//    .x(16),
//    .d(m_dec[3]),
//    .result(decom_out[3])
//);

//decompress_module decompress_inst4 (
//    .x(16),
//    .d(m_dec[4]),
//    .result(decom_out[4])
//);

//decompress_module decompress_inst5 (
//    .x(16),
//    .d(m_dec[5]),
//    .result(decom_out[5])
//);

//decompress_module decompress_inst6 (
//    .x(16),
//    .d(m_dec[6]),
//    .result(decom_out[6])
//);

//decompress_module decompress_inst7 (
//    .x(16),
//    .d(m_dec[7]),
//    .result(decom_out[7])
//);

//decompress_module decompress_inst8 (
//    .x(16),
//    .d(m_dec[8]),
//    .result(decom_out[8])
//);

//decompress_module decompress_inst9 (
//    .x(16),
//    .d(m_dec[9]),
//    .result(decom_out[9])
//);

//decompress_module decompress_inst10 (
//    .x(16),
//    .d(m_dec[10]),
//    .result(decom_out[10])
//);

//decompress_module decompress_inst11 (
//    .x(16),
//    .d(m_dec[11]),
//    .result(decom_out[11])
//);

//decompress_module decompress_inst12 (
//    .x(16),
//    .d(m_dec[12]),
//    .result(decom_out[12])
//);

//decompress_module decompress_inst13 (
//    .x(16),
//    .d(m_dec[13]),
//    .result(decom_out[13])
//);

//decompress_module decompress_inst14 (
//    .x(16),
//    .d(m_dec[14]),
//    .result(decom_out[14])
//);

//decompress_module decompress_inst15 (
//    .x(16),
//    .d(m_dec[15]),
//    .result(decom_out[15])
//);

//decompress_module decompress_inst16 (
//    .x(16),
//    .d(m_dec[16]),
//    .result(decom_out[16])
//);

//decompress_module decompress_inst17 (
//    .x(16),
//    .d(m_dec[17]),
//    .result(decom_out[17])
//);

//decompress_module decompress_inst18 (
//    .x(16),
//    .d(m_dec[18]),
//    .result(decom_out[18])
//);

//decompress_module decompress_inst19 (
//    .x(16),
//    .d(m_dec[19]),
//    .result(decom_out[19])
//);

//decompress_module decompress_inst20 (
//    .x(16),
//    .d(m_dec[20]),
//    .result(decom_out[20])
//);

//decompress_module decompress_inst21 (
//    .x(16),
//    .d(m_dec[21]),
//    .result(decom_out[21])
//);

//decompress_module decompress_inst22 (
//    .x(16),
//    .d(m_dec[22]),
//    .result(decom_out[22])
//);

//decompress_module decompress_inst23 (
//    .x(16),
//    .d(m_dec[23]),
//    .result(decom_out[23])
//);

//decompress_module decompress_inst24 (
//    .x(16),
//    .d(m_dec[24]),
//    .result(decom_out[24])
//);

//decompress_module decompress_inst25 (
//    .x(16),
//    .d(m_dec[25]),
//    .result(decom_out[25])
//);

//decompress_module decompress_inst26 (
//    .x(16),
//    .d(m_dec[26]),
//    .result(decom_out[26])
//);

//decompress_module decompress_inst27 (
//    .x(16),
//    .d(m_dec[27]),
//    .result(decom_out[27])
//);

//decompress_module decompress_inst28 (
//    .x(16),
//    .d(m_dec[28]),
//    .result(decom_out[28])
//);

//decompress_module decompress_inst29 (
//    .x(16),
//    .d(m_dec[29]),
//    .result(decom_out[29])
//);

//decompress_module decompress_inst30 (
//    .x(16),
//    .d(m_dec[30]),
//    .result(decom_out[30])
//);

//decompress_module decompress_inst31 (
//    .x(16),
//    .d(m_dec[31]),
//    .result(decom_out[31])
//);

//decompress_module decompress_inst32 (
//    .x(16),
//    .d(m_dec[32]),
//    .result(decom_out[32])
//);

//decompress_module decompress_inst33 (
//    .x(16),
//    .d(m_dec[33]),
//    .result(decom_out[33])
//);

//decompress_module decompress_inst34 (
//    .x(16),
//    .d(m_dec[34]),
//    .result(decom_out[34])
//);

//decompress_module decompress_inst35 (
//    .x(16),
//    .d(m_dec[35]),
//    .result(decom_out[35])
//);

//decompress_module decompress_inst36 (
//    .x(16),
//    .d(m_dec[36]),
//    .result(decom_out[36])
//);

//decompress_module decompress_inst37 (
//    .x(16),
//    .d(m_dec[37]),
//    .result(decom_out[37])
//);

//decompress_module decompress_inst38 (
//    .x(16),
//    .d(m_dec[38]),
//    .result(decom_out[38])
//);

//decompress_module decompress_inst39 (
//    .x(16),
//    .d(m_dec[39]),
//    .result(decom_out[39])
//);

//decompress_module decompress_inst40 (
//    .x(16),
//    .d(m_dec[40]),
//    .result(decom_out[40])
//);

//decompress_module decompress_inst41 (
//    .x(16),
//    .d(m_dec[41]),
//    .result(decom_out[41])
//);

//decompress_module decompress_inst42 (
//    .x(16),
//    .d(m_dec[42]),
//    .result(decom_out[42])
//);

//decompress_module decompress_inst43 (
//    .x(16),
//    .d(m_dec[43]),
//    .result(decom_out[43])
//);

//decompress_module decompress_inst44 (
//    .x(16),
//    .d(m_dec[44]),
//    .result(decom_out[44])
//);

//decompress_module decompress_inst45 (
//    .x(16),
//    .d(m_dec[45]),
//    .result(decom_out[45])
//);

//decompress_module decompress_inst46 (
//    .x(16),
//    .d(m_dec[46]),
//    .result(decom_out[46])
//);

//decompress_module decompress_inst47 (
//    .x(16),
//    .d(m_dec[47]),
//    .result(decom_out[47])
//);

//decompress_module decompress_inst48 (
//    .x(16),
//    .d(m_dec[48]),
//    .result(decom_out[48])
//);

//decompress_module decompress_inst49 (
//    .x(16),
//    .d(m_dec[49]),
//    .result(decom_out[49])
//);

//decompress_module decompress_inst50 (
//    .x(16),
//    .d(m_dec[50]),
//    .result(decom_out[50])
//);

//decompress_module decompress_inst51 (
//    .x(16),
//    .d(m_dec[51]),
//    .result(decom_out[51])
//);

//decompress_module decompress_inst52 (
//    .x(16),
//    .d(m_dec[52]),
//    .result(decom_out[52])
//);

//decompress_module decompress_inst53 (
//    .x(16),
//    .d(m_dec[53]),
//    .result(decom_out[53])
//);

//decompress_module decompress_inst54 (
//    .x(16),
//    .d(m_dec[54]),
//    .result(decom_out[54])
//);

//decompress_module decompress_inst55 (
//    .x(16),
//    .d(m_dec[55]),
//    .result(decom_out[55])
//);

//decompress_module decompress_inst56 (
//    .x(16),
//    .d(m_dec[56]),
//    .result(decom_out[56])
//);

//decompress_module decompress_inst57 (
//    .x(16),
//    .d(m_dec[57]),
//    .result(decom_out[57])
//);

//decompress_module decompress_inst58 (
//    .x(16),
//    .d(m_dec[58]),
//    .result(decom_out[58])
//);

//decompress_module decompress_inst59 (
//    .x(16),
//    .d(m_dec[59]),
//    .result(decom_out[59])
//);

//decompress_module decompress_inst60 (
//    .x(16),
//    .d(m_dec[60]),
//    .result(decom_out[60])
//);

//decompress_module decompress_inst61 (
//    .x(16),
//    .d(m_dec[61]),
//    .result(decom_out[61])
//);

//decompress_module decompress_inst62 (
//    .x(16),
//    .d(m_dec[62]),
//    .result(decom_out[62])
//);

//decompress_module decompress_inst63 (
//    .x(16),
//    .d(m_dec[63]),
//    .result(decom_out[63])
//);

//decompress_module decompress_inst64 (
//    .x(16),
//    .d(m_dec[64]),
//    .result(decom_out[64])
//);

//decompress_module decompress_inst65 (
//    .x(16),
//    .d(m_dec[65]),
//    .result(decom_out[65])
//);

//decompress_module decompress_inst66 (
//    .x(16),
//    .d(m_dec[66]),
//    .result(decom_out[66])
//);

//decompress_module decompress_inst67 (
//    .x(16),
//    .d(m_dec[67]),
//    .result(decom_out[67])
//);

//decompress_module decompress_inst68 (
//    .x(16),
//    .d(m_dec[68]),
//    .result(decom_out[68])
//);

//decompress_module decompress_inst69 (
//    .x(16),
//    .d(m_dec[69]),
//    .result(decom_out[69])
//);

//decompress_module decompress_inst70 (
//    .x(16),
//    .d(m_dec[70]),
//    .result(decom_out[70])
//);

//decompress_module decompress_inst71 (
//    .x(16),
//    .d(m_dec[71]),
//    .result(decom_out[71])
//);

//decompress_module decompress_inst72 (
//    .x(16),
//    .d(m_dec[72]),
//    .result(decom_out[72])
//);

//decompress_module decompress_inst73 (
//    .x(16),
//    .d(m_dec[73]),
//    .result(decom_out[73])
//);

//decompress_module decompress_inst74 (
//    .x(16),
//    .d(m_dec[74]),
//    .result(decom_out[74])
//);

//decompress_module decompress_inst75 (
//    .x(16),
//    .d(m_dec[75]),
//    .result(decom_out[75])
//);

//decompress_module decompress_inst76 (
//    .x(16),
//    .d(m_dec[76]),
//    .result(decom_out[76])
//);

//decompress_module decompress_inst77 (
//    .x(16),
//    .d(m_dec[77]),
//    .result(decom_out[77])
//);

//decompress_module decompress_inst78 (
//    .x(16),
//    .d(m_dec[78]),
//    .result(decom_out[78])
//);

//decompress_module decompress_inst79 (
//    .x(16),
//    .d(m_dec[79]),
//    .result(decom_out[79])
//);

//decompress_module decompress_inst80 (
//    .x(16),
//    .d(m_dec[80]),
//    .result(decom_out[80])
//);

//decompress_module decompress_inst81 (
//    .x(16),
//    .d(m_dec[81]),
//    .result(decom_out[81])
//);

//decompress_module decompress_inst82 (
//    .x(16),
//    .d(m_dec[82]),
//    .result(decom_out[82])
//);

//decompress_module decompress_inst83 (
//    .x(16),
//    .d(m_dec[83]),
//    .result(decom_out[83])
//);

//decompress_module decompress_inst84 (
//    .x(16),
//    .d(m_dec[84]),
//    .result(decom_out[84])
//);

//decompress_module decompress_inst85 (
//    .x(16),
//    .d(m_dec[85]),
//    .result(decom_out[85])
//);

//decompress_module decompress_inst86 (
//    .x(16),
//    .d(m_dec[86]),
//    .result(decom_out[86])
//);

//decompress_module decompress_inst87 (
//    .x(16),
//    .d(m_dec[87]),
//    .result(decom_out[87])
//);

//decompress_module decompress_inst88 (
//    .x(16),
//    .d(m_dec[88]),
//    .result(decom_out[88])
//);

//decompress_module decompress_inst89 (
//    .x(16),
//    .d(m_dec[89]),
//    .result(decom_out[89])
//);

//decompress_module decompress_inst90 (
//    .x(16),
//    .d(m_dec[90]),
//    .result(decom_out[90])
//);

//decompress_module decompress_inst91 (
//    .x(16),
//    .d(m_dec[91]),
//    .result(decom_out[91])
//);

//decompress_module decompress_inst92 (
//    .x(16),
//    .d(m_dec[92]),
//    .result(decom_out[92])
//);

//decompress_module decompress_inst93 (
//    .x(16),
//    .d(m_dec[93]),
//    .result(decom_out[93])
//);

//decompress_module decompress_inst94 (
//    .x(16),
//    .d(m_dec[94]),
//    .result(decom_out[94])
//);

//decompress_module decompress_inst95 (
//    .x(16),
//    .d(m_dec[95]),
//    .result(decom_out[95])
//);

//decompress_module decompress_inst96 (
//    .x(16),
//    .d(m_dec[96]),
//    .result(decom_out[96])
//);

//decompress_module decompress_inst97 (
//    .x(16),
//    .d(m_dec[97]),
//    .result(decom_out[97])
//);

//decompress_module decompress_inst98 (
//    .x(16),
//    .d(m_dec[98]),
//    .result(decom_out[98])
//);

//decompress_module decompress_inst99 (
//    .x(16),
//    .d(m_dec[99]),
//    .result(decom_out[99])
//);

//decompress_module decompress_inst100 (
//    .x(16),
//    .d(m_dec[100]),
//    .result(decom_out[100])
//);

//decompress_module decompress_inst101 (
//    .x(16),
//    .d(m_dec[101]),
//    .result(decom_out[101])
//);

//decompress_module decompress_inst102 (
//    .x(16),
//    .d(m_dec[102]),
//    .result(decom_out[102])
//);

//decompress_module decompress_inst103 (
//    .x(16),
//    .d(m_dec[103]),
//    .result(decom_out[103])
//);

//decompress_module decompress_inst104 (
//    .x(16),
//    .d(m_dec[104]),
//    .result(decom_out[104])
//);

//decompress_module decompress_inst105 (
//    .x(16),
//    .d(m_dec[105]),
//    .result(decom_out[105])
//);

//decompress_module decompress_inst106 (
//    .x(16),
//    .d(m_dec[106]),
//    .result(decom_out[106])
//);

//decompress_module decompress_inst107 (
//    .x(16),
//    .d(m_dec[107]),
//    .result(decom_out[107])
//);

//decompress_module decompress_inst108 (
//    .x(16),
//    .d(m_dec[108]),
//    .result(decom_out[108])
//);

//decompress_module decompress_inst109 (
//    .x(16),
//    .d(m_dec[109]),
//    .result(decom_out[109])
//);

//decompress_module decompress_inst110 (
//    .x(16),
//    .d(m_dec[110]),
//    .result(decom_out[110])
//);

//decompress_module decompress_inst111 (
//    .x(16),
//    .d(m_dec[111]),
//    .result(decom_out[111])
//);

//decompress_module decompress_inst112 (
//    .x(16),
//    .d(m_dec[112]),
//    .result(decom_out[112])
//);

//decompress_module decompress_inst113 (
//    .x(16),
//    .d(m_dec[113]),
//    .result(decom_out[113])
//);

//decompress_module decompress_inst114 (
//    .x(16),
//    .d(m_dec[114]),
//    .result(decom_out[114])
//);

//decompress_module decompress_inst115 (
//    .x(16),
//    .d(m_dec[115]),
//    .result(decom_out[115])
//);

//decompress_module decompress_inst116 (
//    .x(16),
//    .d(m_dec[116]),
//    .result(decom_out[116])
//);

//decompress_module decompress_inst117 (
//    .x(16),
//    .d(m_dec[117]),
//    .result(decom_out[117])
//);

//decompress_module decompress_inst118 (
//    .x(16),
//    .d(m_dec[118]),
//    .result(decom_out[118])
//);

//decompress_module decompress_inst119 (
//    .x(16),
//    .d(m_dec[119]),
//    .result(decom_out[119])
//);

//decompress_module decompress_inst120 (
//    .x(16),
//    .d(m_dec[120]),
//    .result(decom_out[120])
//);

//decompress_module decompress_inst121 (
//    .x(16),
//    .d(m_dec[121]),
//    .result(decom_out[121])
//);

//decompress_module decompress_inst122 (
//    .x(16),
//    .d(m_dec[122]),
//    .result(decom_out[122])
//);

//decompress_module decompress_inst123 (
//    .x(16),
//    .d(m_dec[123]),
//    .result(decom_out[123])
//);

//decompress_module decompress_inst124 (
//    .x(16),
//    .d(m_dec[124]),
//    .result(decom_out[124])
//);

//decompress_module decompress_inst125 (
//    .x(16),
//    .d(m_dec[125]),
//    .result(decom_out[125])
//);

//decompress_module decompress_inst126 (
//    .x(16),
//    .d(m_dec[126]),
//    .result(decom_out[126])
//);

//decompress_module decompress_inst127 (
//    .x(16),
//    .d(m_dec[127]),
//    .result(decom_out[127])
//);

//decompress_module decompress_inst128 (
//    .x(16),
//    .d(m_dec[128]),
//    .result(decom_out[128])
//);

//decompress_module decompress_inst129 (
//    .x(16),
//    .d(m_dec[129]),
//    .result(decom_out[129])
//);

//decompress_module decompress_inst130 (
//    .x(16),
//    .d(m_dec[130]),
//    .result(decom_out[130])
//);

//decompress_module decompress_inst131 (
//    .x(16),
//    .d(m_dec[131]),
//    .result(decom_out[131])
//);

//decompress_module decompress_inst132 (
//    .x(16),
//    .d(m_dec[132]),
//    .result(decom_out[132])
//);

//decompress_module decompress_inst133 (
//    .x(16),
//    .d(m_dec[133]),
//    .result(decom_out[133])
//);

//decompress_module decompress_inst134 (
//    .x(16),
//    .d(m_dec[134]),
//    .result(decom_out[134])
//);

//decompress_module decompress_inst135 (
//    .x(16),
//    .d(m_dec[135]),
//    .result(decom_out[135])
//);

//decompress_module decompress_inst136 (
//    .x(16),
//    .d(m_dec[136]),
//    .result(decom_out[136])
//);

//decompress_module decompress_inst137 (
//    .x(16),
//    .d(m_dec[137]),
//    .result(decom_out[137])
//);

//decompress_module decompress_inst138 (
//    .x(16),
//    .d(m_dec[138]),
//    .result(decom_out[138])
//);

//decompress_module decompress_inst139 (
//    .x(16),
//    .d(m_dec[139]),
//    .result(decom_out[139])
//);

//decompress_module decompress_inst140 (
//    .x(16),
//    .d(m_dec[140]),
//    .result(decom_out[140])
//);

//decompress_module decompress_inst141 (
//    .x(16),
//    .d(m_dec[141]),
//    .result(decom_out[141])
//);

//decompress_module decompress_inst142 (
//    .x(16),
//    .d(m_dec[142]),
//    .result(decom_out[142])
//);

//decompress_module decompress_inst143 (
//    .x(16),
//    .d(m_dec[143]),
//    .result(decom_out[143])
//);

//decompress_module decompress_inst144 (
//    .x(16),
//    .d(m_dec[144]),
//    .result(decom_out[144])
//);

//decompress_module decompress_inst145 (
//    .x(16),
//    .d(m_dec[145]),
//    .result(decom_out[145])
//);

//decompress_module decompress_inst146 (
//    .x(16),
//    .d(m_dec[146]),
//    .result(decom_out[146])
//);

//decompress_module decompress_inst147 (
//    .x(16),
//    .d(m_dec[147]),
//    .result(decom_out[147])
//);

//decompress_module decompress_inst148 (
//    .x(16),
//    .d(m_dec[148]),
//    .result(decom_out[148])
//);

//decompress_module decompress_inst149 (
//    .x(16),
//    .d(m_dec[149]),
//    .result(decom_out[149])
//);

//decompress_module decompress_inst150 (
//    .x(16),
//    .d(m_dec[150]),
//    .result(decom_out[150])
//);

//decompress_module decompress_inst151 (
//    .x(16),
//    .d(m_dec[151]),
//    .result(decom_out[151])
//);

//decompress_module decompress_inst152 (
//    .x(16),
//    .d(m_dec[152]),
//    .result(decom_out[152])
//);

//decompress_module decompress_inst153 (
//    .x(16),
//    .d(m_dec[153]),
//    .result(decom_out[153])
//);

//decompress_module decompress_inst154 (
//    .x(16),
//    .d(m_dec[154]),
//    .result(decom_out[154])
//);

//decompress_module decompress_inst155 (
//    .x(16),
//    .d(m_dec[155]),
//    .result(decom_out[155])
//);

//decompress_module decompress_inst156 (
//    .x(16),
//    .d(m_dec[156]),
//    .result(decom_out[156])
//);

//decompress_module decompress_inst157 (
//    .x(16),
//    .d(m_dec[157]),
//    .result(decom_out[157])
//);

//decompress_module decompress_inst158 (
//    .x(16),
//    .d(m_dec[158]),
//    .result(decom_out[158])
//);

//decompress_module decompress_inst159 (
//    .x(16),
//    .d(m_dec[159]),
//    .result(decom_out[159])
//);

//decompress_module decompress_inst160 (
//    .x(16),
//    .d(m_dec[160]),
//    .result(decom_out[160])
//);

//decompress_module decompress_inst161 (
//    .x(16),
//    .d(m_dec[161]),
//    .result(decom_out[161])
//);

//decompress_module decompress_inst162 (
//    .x(16),
//    .d(m_dec[162]),
//    .result(decom_out[162])
//);

//decompress_module decompress_inst163 (
//    .x(16),
//    .d(m_dec[163]),
//    .result(decom_out[163])
//);

//decompress_module decompress_inst164 (
//    .x(16),
//    .d(m_dec[164]),
//    .result(decom_out[164])
//);

//decompress_module decompress_inst165 (
//    .x(16),
//    .d(m_dec[165]),
//    .result(decom_out[165])
//);

//decompress_module decompress_inst166 (
//    .x(16),
//    .d(m_dec[166]),
//    .result(decom_out[166])
//);

//decompress_module decompress_inst167 (
//    .x(16),
//    .d(m_dec[167]),
//    .result(decom_out[167])
//);

//decompress_module decompress_inst168 (
//    .x(16),
//    .d(m_dec[168]),
//    .result(decom_out[168])
//);

//decompress_module decompress_inst169 (
//    .x(16),
//    .d(m_dec[169]),
//    .result(decom_out[169])
//);

//decompress_module decompress_inst170 (
//    .x(16),
//    .d(m_dec[170]),
//    .result(decom_out[170])
//);

//decompress_module decompress_inst171 (
//    .x(16),
//    .d(m_dec[171]),
//    .result(decom_out[171])
//);

//decompress_module decompress_inst172 (
//    .x(16),
//    .d(m_dec[172]),
//    .result(decom_out[172])
//);

//decompress_module decompress_inst173 (
//    .x(16),
//    .d(m_dec[173]),
//    .result(decom_out[173])
//);

//decompress_module decompress_inst174 (
//    .x(16),
//    .d(m_dec[174]),
//    .result(decom_out[174])
//);

//decompress_module decompress_inst175 (
//    .x(16),
//    .d(m_dec[175]),
//    .result(decom_out[175])
//);

//decompress_module decompress_inst176 (
//    .x(16),
//    .d(m_dec[176]),
//    .result(decom_out[176])
//);

//decompress_module decompress_inst177 (
//    .x(16),
//    .d(m_dec[177]),
//    .result(decom_out[177])
//);

//decompress_module decompress_inst178 (
//    .x(16),
//    .d(m_dec[178]),
//    .result(decom_out[178])
//);

//decompress_module decompress_inst179 (
//    .x(16),
//    .d(m_dec[179]),
//    .result(decom_out[179])
//);

//decompress_module decompress_inst180 (
//    .x(16),
//    .d(m_dec[180]),
//    .result(decom_out[180])
//);

//decompress_module decompress_inst181 (
//    .x(16),
//    .d(m_dec[181]),
//    .result(decom_out[181])
//);

//decompress_module decompress_inst182 (
//    .x(16),
//    .d(m_dec[182]),
//    .result(decom_out[182])
//);

//decompress_module decompress_inst183 (
//    .x(16),
//    .d(m_dec[183]),
//    .result(decom_out[183])
//);

//decompress_module decompress_inst184 (
//    .x(16),
//    .d(m_dec[184]),
//    .result(decom_out[184])
//);

//decompress_module decompress_inst185 (
//    .x(16),
//    .d(m_dec[185]),
//    .result(decom_out[185])
//);

//decompress_module decompress_inst186 (
//    .x(16),
//    .d(m_dec[186]),
//    .result(decom_out[186])
//);

//decompress_module decompress_inst187 (
//    .x(16),
//    .d(m_dec[187]),
//    .result(decom_out[187])
//);

//decompress_module decompress_inst188 (
//    .x(16),
//    .d(m_dec[188]),
//    .result(decom_out[188])
//);

//decompress_module decompress_inst189 (
//    .x(16),
//    .d(m_dec[189]),
//    .result(decom_out[189])
//);

//decompress_module decompress_inst190 (
//    .x(16),
//    .d(m_dec[190]),
//    .result(decom_out[190])
//);

//decompress_module decompress_inst191 (
//    .x(16),
//    .d(m_dec[191]),
//    .result(decom_out[191])
//);

//decompress_module decompress_inst192 (
//    .x(16),
//    .d(m_dec[192]),
//    .result(decom_out[192])
//);

//decompress_module decompress_inst193 (
//    .x(16),
//    .d(m_dec[193]),
//    .result(decom_out[193])
//);

//decompress_module decompress_inst194 (
//    .x(16),
//    .d(m_dec[194]),
//    .result(decom_out[194])
//);

//decompress_module decompress_inst195 (
//    .x(16),
//    .d(m_dec[195]),
//    .result(decom_out[195])
//);

//decompress_module decompress_inst196 (
//    .x(16),
//    .d(m_dec[196]),
//    .result(decom_out[196])
//);

//decompress_module decompress_inst197 (
//    .x(16),
//    .d(m_dec[197]),
//    .result(decom_out[197])
//);

//decompress_module decompress_inst198 (
//    .x(16),
//    .d(m_dec[198]),
//    .result(decom_out[198])
//);

//decompress_module decompress_inst199 (
//    .x(16),
//    .d(m_dec[199]),
//    .result(decom_out[199])
//);

//decompress_module decompress_inst200 (
//    .x(16),
//    .d(m_dec[200]),
//    .result(decom_out[200])
//);

//decompress_module decompress_inst201 (
//    .x(16),
//    .d(m_dec[201]),
//    .result(decom_out[201])
//);

//decompress_module decompress_inst202 (
//    .x(16),
//    .d(m_dec[202]),
//    .result(decom_out[202])
//);

//decompress_module decompress_inst203 (
//    .x(16),
//    .d(m_dec[203]),
//    .result(decom_out[203])
//);

//decompress_module decompress_inst204 (
//    .x(16),
//    .d(m_dec[204]),
//    .result(decom_out[204])
//);

//decompress_module decompress_inst205 (
//    .x(16),
//    .d(m_dec[205]),
//    .result(decom_out[205])
//);

//decompress_module decompress_inst206 (
//    .x(16),
//    .d(m_dec[206]),
//    .result(decom_out[206])
//);

//decompress_module decompress_inst207 (
//    .x(16),
//    .d(m_dec[207]),
//    .result(decom_out[207])
//);

//decompress_module decompress_inst208 (
//    .x(16),
//    .d(m_dec[208]),
//    .result(decom_out[208])
//);

//decompress_module decompress_inst209 (
//    .x(16),
//    .d(m_dec[209]),
//    .result(decom_out[209])
//);

//decompress_module decompress_inst210 (
//    .x(16),
//    .d(m_dec[210]),
//    .result(decom_out[210])
//);

//decompress_module decompress_inst211 (
//    .x(16),
//    .d(m_dec[211]),
//    .result(decom_out[211])
//);

//decompress_module decompress_inst212 (
//    .x(16),
//    .d(m_dec[212]),
//    .result(decom_out[212])
//);

//decompress_module decompress_inst213 (
//    .x(16),
//    .d(m_dec[213]),
//    .result(decom_out[213])
//);

//decompress_module decompress_inst214 (
//    .x(16),
//    .d(m_dec[214]),
//    .result(decom_out[214])
//);

//decompress_module decompress_inst215 (
//    .x(16),
//    .d(m_dec[215]),
//    .result(decom_out[215])
//);

//decompress_module decompress_inst216 (
//    .x(16),
//    .d(m_dec[216]),
//    .result(decom_out[216])
//);

//decompress_module decompress_inst217 (
//    .x(16),
//    .d(m_dec[217]),
//    .result(decom_out[217])
//);

//decompress_module decompress_inst218 (
//    .x(16),
//    .d(m_dec[218]),
//    .result(decom_out[218])
//);

//decompress_module decompress_inst219 (
//    .x(16),
//    .d(m_dec[219]),
//    .result(decom_out[219])
//);

//decompress_module decompress_inst220 (
//    .x(16),
//    .d(m_dec[220]),
//    .result(decom_out[220])
//);

//decompress_module decompress_inst221 (
//    .x(16),
//    .d(m_dec[221]),
//    .result(decom_out[221])
//);

//decompress_module decompress_inst222 (
//    .x(16),
//    .d(m_dec[222]),
//    .result(decom_out[222])
//);

//decompress_module decompress_inst223 (
//    .x(16),
//    .d(m_dec[223]),
//    .result(decom_out[223])
//);

//decompress_module decompress_inst224 (
//    .x(16),
//    .d(m_dec[224]),
//    .result(decom_out[224])
//);

//decompress_module decompress_inst225 (
//    .x(16),
//    .d(m_dec[225]),
//    .result(decom_out[225])
//);

//decompress_module decompress_inst226 (
//    .x(16),
//    .d(m_dec[226]),
//    .result(decom_out[226])
//);

//decompress_module decompress_inst227 (
//    .x(16),
//    .d(m_dec[227]),
//    .result(decom_out[227])
//);

//decompress_module decompress_inst228 (
//    .x(16),
//    .d(m_dec[228]),
//    .result(decom_out[228])
//);

//decompress_module decompress_inst229 (
//    .x(16),
//    .d(m_dec[229]),
//    .result(decom_out[229])
//);

//decompress_module decompress_inst230 (
//    .x(16),
//    .d(m_dec[230]),
//    .result(decom_out[230])
//);

//decompress_module decompress_inst231 (
//    .x(16),
//    .d(m_dec[231]),
//    .result(decom_out[231])
//);

//decompress_module decompress_inst232 (
//    .x(16),
//    .d(m_dec[232]),
//    .result(decom_out[232])
//);

//decompress_module decompress_inst233 (
//    .x(16),
//    .d(m_dec[233]),
//    .result(decom_out[233])
//);

//decompress_module decompress_inst234 (
//    .x(16),
//    .d(m_dec[234]),
//    .result(decom_out[234])
//);

//decompress_module decompress_inst235 (
//    .x(16),
//    .d(m_dec[235]),
//    .result(decom_out[235])
//);

//decompress_module decompress_inst236 (
//    .x(16),
//    .d(m_dec[236]),
//    .result(decom_out[236])
//);

//decompress_module decompress_inst237 (
//    .x(16),
//    .d(m_dec[237]),
//    .result(decom_out[237])
//);

//decompress_module decompress_inst238 (
//    .x(16),
//    .d(m_dec[238]),
//    .result(decom_out[238])
//);

//decompress_module decompress_inst239 (
//    .x(16),
//    .d(m_dec[239]),
//    .result(decom_out[239])
//);

//decompress_module decompress_inst240 (
//    .x(16),
//    .d(m_dec[240]),
//    .result(decom_out[240])
//);

//decompress_module decompress_inst241 (
//    .x(16),
//    .d(m_dec[241]),
//    .result(decom_out[241])
//);

//decompress_module decompress_inst242 (
//    .x(16),
//    .d(m_dec[242]),
//    .result(decom_out[242])
//);

//decompress_module decompress_inst243 (
//    .x(16),
//    .d(m_dec[243]),
//    .result(decom_out[243])
//);

//decompress_module decompress_inst244 (
//    .x(16),
//    .d(m_dec[244]),
//    .result(decom_out[244])
//);

//decompress_module decompress_inst245 (
//    .x(16),
//    .d(m_dec[245]),
//    .result(decom_out[245])
//);

//decompress_module decompress_inst246 (
//    .x(16),
//    .d(m_dec[246]),
//    .result(decom_out[246])
//);

//decompress_module decompress_inst247 (
//    .x(16),
//    .d(m_dec[247]),
//    .result(decom_out[247])
//);

//decompress_module decompress_inst248 (
//    .x(16),
//    .d(m_dec[248]),
//    .result(decom_out[248])
//);

//decompress_module decompress_inst249 (
//    .x(16),
//    .d(m_dec[249]),
//    .result(decom_out[249])
//);

//decompress_module decompress_inst250 (
//    .x(16),
//    .d(m_dec[250]),
//    .result(decom_out[250])
//);

//decompress_module decompress_inst251 (
//    .x(16),
//    .d(m_dec[251]),
//    .result(decom_out[251])
//);

//decompress_module decompress_inst252 (
//    .x(16),
//    .d(m_dec[252]),
//    .result(decom_out[252])
//);

//decompress_module decompress_inst253 (
//    .x(16),
//    .d(m_dec[253]),
//    .result(decom_out[253])
//);

//decompress_module decompress_inst254 (
//    .x(16),
//    .d(m_dec[254]),
//    .result(decom_out[254])
//);

//decompress_module decompress_inst255 (
//    .x(16),
//    .d(m_dec[255]),
//    .result(decom_out[255])
//);
////v = NTT_inverse(T_hat x Y) + e2 + u

//assign e2_ext[0] = {30'd0, e2[0]};
//assign e2_ext[1] = {30'd0, e2[1]};
//assign e2_ext[2] = {30'd0, e2[2]};
//assign e2_ext[3] = {30'd0, e2[3]};
//assign e2_ext[4] = {30'd0, e2[4]};
//assign e2_ext[5] = {30'd0, e2[5]};
//assign e2_ext[6] = {30'd0, e2[6]};
//assign e2_ext[7] = {30'd0, e2[7]};
//assign e2_ext[8] = {30'd0, e2[8]};
//assign e2_ext[9] = {30'd0, e2[9]};
//assign e2_ext[10] = {30'd0, e2[10]};
//assign e2_ext[11] = {30'd0, e2[11]};
//assign e2_ext[12] = {30'd0, e2[12]};
//assign e2_ext[13] = {30'd0, e2[13]};
//assign e2_ext[14] = {30'd0, e2[14]};
//assign e2_ext[15] = {30'd0, e2[15]};
//assign e2_ext[16] = {30'd0, e2[16]};
//assign e2_ext[17] = {30'd0, e2[17]};
//assign e2_ext[18] = {30'd0, e2[18]};
//assign e2_ext[19] = {30'd0, e2[19]};
//assign e2_ext[20] = {30'd0, e2[20]};
//assign e2_ext[21] = {30'd0, e2[21]};
//assign e2_ext[22] = {30'd0, e2[22]};
//assign e2_ext[23] = {30'd0, e2[23]};
//assign e2_ext[24] = {30'd0, e2[24]};
//assign e2_ext[25] = {30'd0, e2[25]};
//assign e2_ext[26] = {30'd0, e2[26]};
//assign e2_ext[27] = {30'd0, e2[27]};
//assign e2_ext[28] = {30'd0, e2[28]};
//assign e2_ext[29] = {30'd0, e2[29]};
//assign e2_ext[30] = {30'd0, e2[30]};
//assign e2_ext[31] = {30'd0, e2[31]};
//assign e2_ext[32] = {30'd0, e2[32]};
//assign e2_ext[33] = {30'd0, e2[33]};
//assign e2_ext[34] = {30'd0, e2[34]};
//assign e2_ext[35] = {30'd0, e2[35]};
//assign e2_ext[36] = {30'd0, e2[36]};
//assign e2_ext[37] = {30'd0, e2[37]};
//assign e2_ext[38] = {30'd0, e2[38]};
//assign e2_ext[39] = {30'd0, e2[39]};
//assign e2_ext[40] = {30'd0, e2[40]};
//assign e2_ext[41] = {30'd0, e2[41]};
//assign e2_ext[42] = {30'd0, e2[42]};
//assign e2_ext[43] = {30'd0, e2[43]};
//assign e2_ext[44] = {30'd0, e2[44]};
//assign e2_ext[45] = {30'd0, e2[45]};
//assign e2_ext[46] = {30'd0, e2[46]};
//assign e2_ext[47] = {30'd0, e2[47]};
//assign e2_ext[48] = {30'd0, e2[48]};
//assign e2_ext[49] = {30'd0, e2[49]};
//assign e2_ext[50] = {30'd0, e2[50]};
//assign e2_ext[51] = {30'd0, e2[51]};
//assign e2_ext[52] = {30'd0, e2[52]};
//assign e2_ext[53] = {30'd0, e2[53]};
//assign e2_ext[54] = {30'd0, e2[54]};
//assign e2_ext[55] = {30'd0, e2[55]};
//assign e2_ext[56] = {30'd0, e2[56]};
//assign e2_ext[57] = {30'd0, e2[57]};
//assign e2_ext[58] = {30'd0, e2[58]};
//assign e2_ext[59] = {30'd0, e2[59]};
//assign e2_ext[60] = {30'd0, e2[60]};
//assign e2_ext[61] = {30'd0, e2[61]};
//assign e2_ext[62] = {30'd0, e2[62]};
//assign e2_ext[63] = {30'd0, e2[63]};
//assign e2_ext[64] = {30'd0, e2[64]};
//assign e2_ext[65] = {30'd0, e2[65]};
//assign e2_ext[66] = {30'd0, e2[66]};
//assign e2_ext[67] = {30'd0, e2[67]};
//assign e2_ext[68] = {30'd0, e2[68]};
//assign e2_ext[69] = {30'd0, e2[69]};
//assign e2_ext[70] = {30'd0, e2[70]};
//assign e2_ext[71] = {30'd0, e2[71]};
//assign e2_ext[72] = {30'd0, e2[72]};
//assign e2_ext[73] = {30'd0, e2[73]};
//assign e2_ext[74] = {30'd0, e2[74]};
//assign e2_ext[75] = {30'd0, e2[75]};
//assign e2_ext[76] = {30'd0, e2[76]};
//assign e2_ext[77] = {30'd0, e2[77]};
//assign e2_ext[78] = {30'd0, e2[78]};
//assign e2_ext[79] = {30'd0, e2[79]};
//assign e2_ext[80] = {30'd0, e2[80]};
//assign e2_ext[81] = {30'd0, e2[81]};
//assign e2_ext[82] = {30'd0, e2[82]};
//assign e2_ext[83] = {30'd0, e2[83]};
//assign e2_ext[84] = {30'd0, e2[84]};
//assign e2_ext[85] = {30'd0, e2[85]};
//assign e2_ext[86] = {30'd0, e2[86]};
//assign e2_ext[87] = {30'd0, e2[87]};
//assign e2_ext[88] = {30'd0, e2[88]};
//assign e2_ext[89] = {30'd0, e2[89]};
//assign e2_ext[90] = {30'd0, e2[90]};
//assign e2_ext[91] = {30'd0, e2[91]};
//assign e2_ext[92] = {30'd0, e2[92]};
//assign e2_ext[93] = {30'd0, e2[93]};
//assign e2_ext[94] = {30'd0, e2[94]};
//assign e2_ext[95] = {30'd0, e2[95]};
//assign e2_ext[96] = {30'd0, e2[96]};
//assign e2_ext[97] = {30'd0, e2[97]};
//assign e2_ext[98] = {30'd0, e2[98]};
//assign e2_ext[99] = {30'd0, e2[99]};
//assign e2_ext[100] = {30'd0, e2[100]};
//assign e2_ext[101] = {30'd0, e2[101]};
//assign e2_ext[102] = {30'd0, e2[102]};
//assign e2_ext[103] = {30'd0, e2[103]};
//assign e2_ext[104] = {30'd0, e2[104]};
//assign e2_ext[105] = {30'd0, e2[105]};
//assign e2_ext[106] = {30'd0, e2[106]};
//assign e2_ext[107] = {30'd0, e2[107]};
//assign e2_ext[108] = {30'd0, e2[108]};
//assign e2_ext[109] = {30'd0, e2[109]};
//assign e2_ext[110] = {30'd0, e2[110]};
//assign e2_ext[111] = {30'd0, e2[111]};
//assign e2_ext[112] = {30'd0, e2[112]};
//assign e2_ext[113] = {30'd0, e2[113]};
//assign e2_ext[114] = {30'd0, e2[114]};
//assign e2_ext[115] = {30'd0, e2[115]};
//assign e2_ext[116] = {30'd0, e2[116]};
//assign e2_ext[117] = {30'd0, e2[117]};
//assign e2_ext[118] = {30'd0, e2[118]};
//assign e2_ext[119] = {30'd0, e2[119]};
//assign e2_ext[120] = {30'd0, e2[120]};
//assign e2_ext[121] = {30'd0, e2[121]};
//assign e2_ext[122] = {30'd0, e2[122]};
//assign e2_ext[123] = {30'd0, e2[123]};
//assign e2_ext[124] = {30'd0, e2[124]};
//assign e2_ext[125] = {30'd0, e2[125]};
//assign e2_ext[126] = {30'd0, e2[126]};
//assign e2_ext[127] = {30'd0, e2[127]};
//assign e2_ext[128] = {30'd0, e2[128]};
//assign e2_ext[129] = {30'd0, e2[129]};
//assign e2_ext[130] = {30'd0, e2[130]};
//assign e2_ext[131] = {30'd0, e2[131]};
//assign e2_ext[132] = {30'd0, e2[132]};
//assign e2_ext[133] = {30'd0, e2[133]};
//assign e2_ext[134] = {30'd0, e2[134]};
//assign e2_ext[135] = {30'd0, e2[135]};
//assign e2_ext[136] = {30'd0, e2[136]};
//assign e2_ext[137] = {30'd0, e2[137]};
//assign e2_ext[138] = {30'd0, e2[138]};
//assign e2_ext[139] = {30'd0, e2[139]};
//assign e2_ext[140] = {30'd0, e2[140]};
//assign e2_ext[141] = {30'd0, e2[141]};
//assign e2_ext[142] = {30'd0, e2[142]};
//assign e2_ext[143] = {30'd0, e2[143]};
//assign e2_ext[144] = {30'd0, e2[144]};
//assign e2_ext[145] = {30'd0, e2[145]};
//assign e2_ext[146] = {30'd0, e2[146]};
//assign e2_ext[147] = {30'd0, e2[147]};
//assign e2_ext[148] = {30'd0, e2[148]};
//assign e2_ext[149] = {30'd0, e2[149]};
//assign e2_ext[150] = {30'd0, e2[150]};
//assign e2_ext[151] = {30'd0, e2[151]};
//assign e2_ext[152] = {30'd0, e2[152]};
//assign e2_ext[153] = {30'd0, e2[153]};
//assign e2_ext[154] = {30'd0, e2[154]};
//assign e2_ext[155] = {30'd0, e2[155]};
//assign e2_ext[156] = {30'd0, e2[156]};
//assign e2_ext[157] = {30'd0, e2[157]};
//assign e2_ext[158] = {30'd0, e2[158]};
//assign e2_ext[159] = {30'd0, e2[159]};
//assign e2_ext[160] = {30'd0, e2[160]};
//assign e2_ext[161] = {30'd0, e2[161]};
//assign e2_ext[162] = {30'd0, e2[162]};
//assign e2_ext[163] = {30'd0, e2[163]};
//assign e2_ext[164] = {30'd0, e2[164]};
//assign e2_ext[165] = {30'd0, e2[165]};
//assign e2_ext[166] = {30'd0, e2[166]};
//assign e2_ext[167] = {30'd0, e2[167]};
//assign e2_ext[168] = {30'd0, e2[168]};
//assign e2_ext[169] = {30'd0, e2[169]};
//assign e2_ext[170] = {30'd0, e2[170]};
//assign e2_ext[171] = {30'd0, e2[171]};
//assign e2_ext[172] = {30'd0, e2[172]};
//assign e2_ext[173] = {30'd0, e2[173]};
//assign e2_ext[174] = {30'd0, e2[174]};
//assign e2_ext[175] = {30'd0, e2[175]};
//assign e2_ext[176] = {30'd0, e2[176]};
//assign e2_ext[177] = {30'd0, e2[177]};
//assign e2_ext[178] = {30'd0, e2[178]};
//assign e2_ext[179] = {30'd0, e2[179]};
//assign e2_ext[180] = {30'd0, e2[180]};
//assign e2_ext[181] = {30'd0, e2[181]};
//assign e2_ext[182] = {30'd0, e2[182]};
//assign e2_ext[183] = {30'd0, e2[183]};
//assign e2_ext[184] = {30'd0, e2[184]};
//assign e2_ext[185] = {30'd0, e2[185]};
//assign e2_ext[186] = {30'd0, e2[186]};
//assign e2_ext[187] = {30'd0, e2[187]};
//assign e2_ext[188] = {30'd0, e2[188]};
//assign e2_ext[189] = {30'd0, e2[189]};
//assign e2_ext[190] = {30'd0, e2[190]};
//assign e2_ext[191] = {30'd0, e2[191]};
//assign e2_ext[192] = {30'd0, e2[192]};
//assign e2_ext[193] = {30'd0, e2[193]};
//assign e2_ext[194] = {30'd0, e2[194]};
//assign e2_ext[195] = {30'd0, e2[195]};
//assign e2_ext[196] = {30'd0, e2[196]};
//assign e2_ext[197] = {30'd0, e2[197]};
//assign e2_ext[198] = {30'd0, e2[198]};
//assign e2_ext[199] = {30'd0, e2[199]};
//assign e2_ext[200] = {30'd0, e2[200]};
//assign e2_ext[201] = {30'd0, e2[201]};
//assign e2_ext[202] = {30'd0, e2[202]};
//assign e2_ext[203] = {30'd0, e2[203]};
//assign e2_ext[204] = {30'd0, e2[204]};
//assign e2_ext[205] = {30'd0, e2[205]};
//assign e2_ext[206] = {30'd0, e2[206]};
//assign e2_ext[207] = {30'd0, e2[207]};
//assign e2_ext[208] = {30'd0, e2[208]};;
//assign e2_ext[209] = {30'd0, e2[209]};
//assign e2_ext[210] = {30'd0, e2[210]};
//assign e2_ext[211] = {30'd0, e2[211]};
//assign e2_ext[212] = {30'd0, e2[212]};
//assign e2_ext[213] = {30'd0, e2[213]};
//assign e2_ext[214] = {30'd0, e2[214]};
//assign e2_ext[215] = {30'd0, e2[215]};
//assign e2_ext[216] = {30'd0, e2[216]};
//assign e2_ext[217] = {30'd0, e2[217]};
//assign e2_ext[218] = {30'd0, e2[218]};
//assign e2_ext[219] = {30'd0, e2[219]};
//assign e2_ext[220] = {30'd0, e2[220]};
//assign e2_ext[221] = {30'd0, e2[221]};
//assign e2_ext[222] = {30'd0, e2[222]};
//assign e2_ext[223] = {30'd0, e2[223]};
//assign e2_ext[224] = {30'd0, e2[224]};
//assign e2_ext[225] = {30'd0, e2[225]};
//assign e2_ext[226] = {30'd0, e2[226]};
//assign e2_ext[227] = {30'd0, e2[227]};
//assign e2_ext[228] = {30'd0, e2[228]};
//assign e2_ext[229] = {30'd0, e2[229]};
//assign e2_ext[230] = {30'd0, e2[230]};
//assign e2_ext[231] = {30'd0, e2[231]};
//assign e2_ext[232] = {30'd0, e2[232]};
//assign e2_ext[233] = {30'd0, e2[233]};
//assign e2_ext[234] = {30'd0, e2[234]};
//assign e2_ext[235] = {30'd0, e2[235]};
//assign e2_ext[236] = {30'd0, e2[236]};
//assign e2_ext[237] = {30'd0, e2[237]};
//assign e2_ext[238] = {30'd0, e2[238]};
//assign e2_ext[239] = {30'd0, e2[239]};
//assign e2_ext[240] = {30'd0, e2[240]};
//assign e2_ext[241] = {30'd0, e2[241]};
//assign e2_ext[242] = {30'd0, e2[242]};
//assign e2_ext[243] = {30'd0, e2[243]};
//assign e2_ext[244] = {30'd0, e2[244]};
//assign e2_ext[245] = {30'd0, e2[245]};
//assign e2_ext[246] = {30'd0, e2[246]};
//assign e2_ext[247] = {30'd0, e2[247]};
//assign e2_ext[248] = {30'd0, e2[248]};
//assign e2_ext[249] = {30'd0, e2[249]};
//assign e2_ext[250] = {30'd0, e2[250]};
//assign e2_ext[251] = {30'd0, e2[251]};
//assign e2_ext[252] = {30'd0, e2[252]};
//assign e2_ext[253] = {30'd0, e2[253]};
//assign e2_ext[254] = {30'd0, e2[254]};
//assign e2_ext[255] = {30'd0, e2[255]};
//assign v_1[0] = {16'd0, decom_out[0] + v_in_1[0] + e2_ext[0]};
//assign v_1[1] = {16'd0, decom_out[1] + v_in_1[1] + e2_ext[1]};
//assign v_1[2] = {16'd0, decom_out[2] + v_in_1[2] + e2_ext[2]};
//assign v_1[3] = {16'd0, decom_out[3] + v_in_1[3] + e2_ext[3]};
//assign v_1[4] = {16'd0, decom_out[4] + v_in_1[4] + e2_ext[4]};
//assign v_1[5] = {16'd0, decom_out[5] + v_in_1[5] + e2_ext[5]};
//assign v_1[6] = {16'd0, decom_out[6] + v_in_1[6] + e2_ext[6]};
//assign v_1[7] = {16'd0, decom_out[7] + v_in_1[7] + e2_ext[7]};
//assign v_1[8] = {16'd0, decom_out[8] + v_in_1[8] + e2_ext[8]};
//assign v_1[9] = {16'd0, decom_out[9] + v_in_1[9] + e2_ext[9]};
//assign v_1[10] = {16'd0, decom_out[10] + v_in_1[10] + e2_ext[10]};
//assign v_1[11] = {16'd0, decom_out[11] + v_in_1[11] + e2_ext[11]};
//assign v_1[12] = {16'd0, decom_out[12] + v_in_1[12] + e2_ext[12]};
//assign v_1[13] = {16'd0, decom_out[13] + v_in_1[13] + e2_ext[13]};
//assign v_1[14] = {16'd0, decom_out[14] + v_in_1[14] + e2_ext[14]};
//assign v_1[15] = {16'd0, decom_out[15] + v_in_1[15] + e2_ext[15]};
//assign v_1[16] = {16'd0, decom_out[16] + v_in_1[16] + e2_ext[16]};
//assign v_1[17] = {16'd0, decom_out[17] + v_in_1[17] + e2_ext[17]};
//assign v_1[18] = {16'd0, decom_out[18] + v_in_1[18] + e2_ext[18]};
//assign v_1[19] = {16'd0, decom_out[19] + v_in_1[19] + e2_ext[19]};
//assign v_1[20] = {16'd0, decom_out[20] + v_in_1[20] + e2_ext[20]};
//assign v_1[21] = {16'd0, decom_out[21] + v_in_1[21] + e2_ext[21]};
//assign v_1[22] = {16'd0, decom_out[22] + v_in_1[22] + e2_ext[22]};
//assign v_1[23] = {16'd0, decom_out[23] + v_in_1[23] + e2_ext[23]};
//assign v_1[24] = {16'd0, decom_out[24] + v_in_1[24] + e2_ext[24]};
//assign v_1[25] = {16'd0, decom_out[25] + v_in_1[25] + e2_ext[25]};
//assign v_1[26] = {16'd0, decom_out[26] + v_in_1[26] + e2_ext[26]};
//assign v_1[27] = {16'd0, decom_out[27] + v_in_1[27] + e2_ext[27]};
//assign v_1[28] = {16'd0, decom_out[28] + v_in_1[28] + e2_ext[28]};
//assign v_1[29] = {16'd0, decom_out[29] + v_in_1[29] + e2_ext[29]};
//assign v_1[30] = {16'd0, decom_out[30] + v_in_1[30] + e2_ext[30]};
//assign v_1[31] = {16'd0, decom_out[31] + v_in_1[31] + e2_ext[31]};
//assign v_1[32] = {16'd0, decom_out[32] + v_in_1[32] + e2_ext[32]};
//assign v_1[33] = {16'd0, decom_out[33] + v_in_1[33] + e2_ext[33]};
//assign v_1[34] = {16'd0, decom_out[34] + v_in_1[34] + e2_ext[34]};
//assign v_1[35] = {16'd0, decom_out[35] + v_in_1[35] + e2_ext[35]};
//assign v_1[36] = {16'd0, decom_out[36] + v_in_1[36] + e2_ext[36]};
//assign v_1[37] = {16'd0, decom_out[37] + v_in_1[37] + e2_ext[37]};
//assign v_1[38] = {16'd0, decom_out[38] + v_in_1[38] + e2_ext[38]};
//assign v_1[39] = {16'd0, decom_out[39] + v_in_1[39] + e2_ext[39]};
//assign v_1[40] = {16'd0, decom_out[40] + v_in_1[40] + e2_ext[40]};
//assign v_1[41] = {16'd0, decom_out[41] + v_in_1[41] + e2_ext[41]};
//assign v_1[42] = {16'd0, decom_out[42] + v_in_1[42] + e2_ext[42]};
//assign v_1[43] = {16'd0, decom_out[43] + v_in_1[43] + e2_ext[43]};
//assign v_1[44] = {16'd0, decom_out[44] + v_in_1[44] + e2_ext[44]};
//assign v_1[45] = {16'd0, decom_out[45] + v_in_1[45] + e2_ext[45]};
//assign v_1[46] = {16'd0, decom_out[46] + v_in_1[46] + e2_ext[46]};
//assign v_1[47] = {16'd0, decom_out[47] + v_in_1[47] + e2_ext[47]};
//assign v_1[48] = {16'd0, decom_out[48] + v_in_1[48] + e2_ext[48]};
//assign v_1[49] = {16'd0, decom_out[49] + v_in_1[49] + e2_ext[49]};
//assign v_1[50] = {16'd0, decom_out[50] + v_in_1[50] + e2_ext[50]};
//assign v_1[51] = {16'd0, decom_out[51] + v_in_1[51] + e2_ext[51]};
//assign v_1[52] = {16'd0, decom_out[52] + v_in_1[52] + e2_ext[52]};
//assign v_1[53] = {16'd0, decom_out[53] + v_in_1[53] + e2_ext[53]};
//assign v_1[54] = {16'd0, decom_out[54] + v_in_1[54] + e2_ext[54]};
//assign v_1[55] = {16'd0, decom_out[55] + v_in_1[55] + e2_ext[55]};
//assign v_1[56] = {16'd0, decom_out[56] + v_in_1[56] + e2_ext[56]};
//assign v_1[57] = {16'd0, decom_out[57] + v_in_1[57] + e2_ext[57]};
//assign v_1[58] = {16'd0, decom_out[58] + v_in_1[58] + e2_ext[58]};
//assign v_1[59] = {16'd0, decom_out[59] + v_in_1[59] + e2_ext[59]};
//assign v_1[60] = {16'd0, decom_out[60] + v_in_1[60] + e2_ext[60]};
//assign v_1[61] = {16'd0, decom_out[61] + v_in_1[61] + e2_ext[61]};
//assign v_1[62] = {16'd0, decom_out[62] + v_in_1[62] + e2_ext[62]};
//assign v_1[63] = {16'd0, decom_out[63] + v_in_1[63] + e2_ext[63]};
//assign v_1[64] = {16'd0, decom_out[64] + v_in_1[64] + e2_ext[64]};
//assign v_1[65] = {16'd0, decom_out[65] + v_in_1[65] + e2_ext[65]};
//assign v_1[66] = {16'd0, decom_out[66] + v_in_1[66] + e2_ext[66]};
//assign v_1[67] = {16'd0, decom_out[67] + v_in_1[67] + e2_ext[67]};
//assign v_1[68] = {16'd0, decom_out[68] + v_in_1[68] + e2_ext[68]};
//assign v_1[69] = {16'd0, decom_out[69] + v_in_1[69] + e2_ext[69]};
//assign v_1[70] = {16'd0, decom_out[70] + v_in_1[70] + e2_ext[70]};
//assign v_1[71] = {16'd0, decom_out[71] + v_in_1[71] + e2_ext[71]};
//assign v_1[72] = {16'd0, decom_out[72] + v_in_1[72] + e2_ext[72]};
//assign v_1[73] = {16'd0, decom_out[73] + v_in_1[73] + e2_ext[73]};
//assign v_1[74] = {16'd0, decom_out[74] + v_in_1[74] + e2_ext[74]};
//assign v_1[75] = {16'd0, decom_out[75] + v_in_1[75] + e2_ext[75]};
//assign v_1[76] = {16'd0, decom_out[76] + v_in_1[76] + e2_ext[76]};
//assign v_1[77] = {16'd0, decom_out[77] + v_in_1[77] + e2_ext[77]};
//assign v_1[78] = {16'd0, decom_out[78] + v_in_1[78] + e2_ext[78]};
//assign v_1[79] = {16'd0, decom_out[79] + v_in_1[79] + e2_ext[79]};
//assign v_1[80] = {16'd0, decom_out[80] + v_in_1[80] + e2_ext[80]};
//assign v_1[81] = {16'd0, decom_out[81] + v_in_1[81] + e2_ext[81]};
//assign v_1[82] = {16'd0, decom_out[82] + v_in_1[82] + e2_ext[82]};
//assign v_1[83] = {16'd0, decom_out[83] + v_in_1[83] + e2_ext[83]};
//assign v_1[84] = {16'd0, decom_out[84] + v_in_1[84] + e2_ext[84]};
//assign v_1[85] = {16'd0, decom_out[85] + v_in_1[85] + e2_ext[85]};
//assign v_1[86] = {16'd0, decom_out[86] + v_in_1[86] + e2_ext[86]};
//assign v_1[87] = {16'd0, decom_out[87] + v_in_1[87] + e2_ext[87]};
//assign v_1[88] = {16'd0, decom_out[88] + v_in_1[88] + e2_ext[88]};
//assign v_1[89] = {16'd0, decom_out[89] + v_in_1[89] + e2_ext[89]};
//assign v_1[90] = {16'd0, decom_out[90] + v_in_1[90] + e2_ext[90]};
//assign v_1[91] = {16'd0, decom_out[91] + v_in_1[91] + e2_ext[91]};
//assign v_1[92] = {16'd0, decom_out[92] + v_in_1[92] + e2_ext[92]};
//assign v_1[93] = {16'd0, decom_out[93] + v_in_1[93] + e2_ext[93]};
//assign v_1[94] = {16'd0, decom_out[94] + v_in_1[94] + e2_ext[94]};
//assign v_1[95] = {16'd0, decom_out[95] + v_in_1[95] + e2_ext[95]};
//assign v_1[96] = {16'd0, decom_out[96] + v_in_1[96] + e2_ext[96]};
//assign v_1[97] = {16'd0, decom_out[97] + v_in_1[97] + e2_ext[97]};
//assign v_1[98] = {16'd0, decom_out[98] + v_in_1[98] + e2_ext[98]};
//assign v_1[99] = {16'd0, decom_out[99] + v_in_1[99] + e2_ext[99]};
//assign v_1[100] = {16'd0, decom_out[100] + v_in_1[100] + e2_ext[100]};
//assign v_1[101] = {16'd0, decom_out[101] + v_in_1[101] + e2_ext[101]};
//assign v_1[102] = {16'd0, decom_out[102] + v_in_1[102] + e2_ext[102]};
//assign v_1[103] = {16'd0, decom_out[103] + v_in_1[103] + e2_ext[103]};
//assign v_1[104] = {16'd0, decom_out[104] + v_in_1[104] + e2_ext[104]};
//assign v_1[105] = {16'd0, decom_out[105] + v_in_1[105] + e2_ext[105]};
//assign v_1[106] = {16'd0, decom_out[106] + v_in_1[106] + e2_ext[106]};
//assign v_1[107] = {16'd0, decom_out[107] + v_in_1[107] + e2_ext[107]};
//assign v_1[108] = {16'd0, decom_out[108] + v_in_1[108] + e2_ext[108]};
//assign v_1[109] = {16'd0, decom_out[109] + v_in_1[109] + e2_ext[109]};
//assign v_1[110] = {16'd0, decom_out[110] + v_in_1[110] + e2_ext[110]};
//assign v_1[111] = {16'd0, decom_out[111] + v_in_1[111] + e2_ext[111]};
//assign v_1[112] = {16'd0, decom_out[112] + v_in_1[112] + e2_ext[112]};
//assign v_1[113] = {16'd0, decom_out[113] + v_in_1[113] + e2_ext[113]};
//assign v_1[114] = {16'd0, decom_out[114] + v_in_1[114] + e2_ext[114]};
//assign v_1[115] = {16'd0, decom_out[115] + v_in_1[115] + e2_ext[115]};
//assign v_1[116] = {16'd0, decom_out[116] + v_in_1[116] + e2_ext[116]};
//assign v_1[117] = {16'd0, decom_out[117] + v_in_1[117] + e2_ext[117]};
//assign v_1[118] = {16'd0, decom_out[118] + v_in_1[118] + e2_ext[118]};
//assign v_1[119] = {16'd0, decom_out[119] + v_in_1[119] + e2_ext[119]};
//assign v_1[120] = {16'd0, decom_out[120] + v_in_1[120] + e2_ext[120]};
//assign v_1[121] = {16'd0, decom_out[121] + v_in_1[121] + e2_ext[121]};
//assign v_1[122] = {16'd0, decom_out[122] + v_in_1[122] + e2_ext[122]};
//assign v_1[123] = {16'd0, decom_out[123] + v_in_1[123] + e2_ext[123]};
//assign v_1[124] = {16'd0, decom_out[124] + v_in_1[124] + e2_ext[124]};
//assign v_1[125] = {16'd0, decom_out[125] + v_in_1[125] + e2_ext[125]};
//assign v_1[126] = {16'd0, decom_out[126] + v_in_1[126] + e2_ext[126]};
//assign v_1[127] = {16'd0, decom_out[127] + v_in_1[127] + e2_ext[127]};
//assign v_1[128] = {16'd0, decom_out[128] + v_in_1[128] + e2_ext[128]};
//assign v_1[129] = {16'd0, decom_out[129] + v_in_1[129] + e2_ext[129]};
//assign v_1[130] = {16'd0, decom_out[130] + v_in_1[130] + e2_ext[130]};
//assign v_1[131] = {16'd0, decom_out[131] + v_in_1[131] + e2_ext[131]};
//assign v_1[132] = {16'd0, decom_out[132] + v_in_1[132] + e2_ext[132]};
//assign v_1[133] = {16'd0, decom_out[133] + v_in_1[133] + e2_ext[133]};
//assign v_1[134] = {16'd0, decom_out[134] + v_in_1[134] + e2_ext[134]};
//assign v_1[135] = {16'd0, decom_out[135] + v_in_1[135] + e2_ext[135]};
//assign v_1[136] = {16'd0, decom_out[136] + v_in_1[136] + e2_ext[136]};
//assign v_1[137] = {16'd0, decom_out[137] + v_in_1[137] + e2_ext[137]};
//assign v_1[138] = {16'd0, decom_out[138] + v_in_1[138] + e2_ext[138]};
//assign v_1[139] = {16'd0, decom_out[139] + v_in_1[139] + e2_ext[139]};
//assign v_1[140] = {16'd0, decom_out[140] + v_in_1[140] + e2_ext[140]};
//assign v_1[141] = {16'd0, decom_out[141] + v_in_1[141] + e2_ext[141]};
//assign v_1[142] = {16'd0, decom_out[142] + v_in_1[142] + e2_ext[142]};
//assign v_1[143] = {16'd0, decom_out[143] + v_in_1[143] + e2_ext[143]};
//assign v_1[144] = {16'd0, decom_out[144] + v_in_1[144] + e2_ext[144]};
//assign v_1[145] = {16'd0, decom_out[145] + v_in_1[145] + e2_ext[145]};
//assign v_1[146] = {16'd0, decom_out[146] + v_in_1[146] + e2_ext[146]};
//assign v_1[147] = {16'd0, decom_out[147] + v_in_1[147] + e2_ext[147]};
//assign v_1[148] = {16'd0, decom_out[148] + v_in_1[148] + e2_ext[148]};
//assign v_1[149] = {16'd0, decom_out[149] + v_in_1[149] + e2_ext[149]};
//assign v_1[150] = {16'd0, decom_out[150] + v_in_1[150] + e2_ext[150]};
//assign v_1[151] = {16'd0, decom_out[151] + v_in_1[151] + e2_ext[151]};
//assign v_1[152] = {16'd0, decom_out[152] + v_in_1[152] + e2_ext[152]};
//assign v_1[153] = {16'd0, decom_out[153] + v_in_1[153] + e2_ext[153]};
//assign v_1[154] = {16'd0, decom_out[154] + v_in_1[154] + e2_ext[154]};
//assign v_1[155] = {16'd0, decom_out[155] + v_in_1[155] + e2_ext[155]};
//assign v_1[156] = {16'd0, decom_out[156] + v_in_1[156] + e2_ext[156]};
//assign v_1[157] = {16'd0, decom_out[157] + v_in_1[157] + e2_ext[157]};
//assign v_1[158] = {16'd0, decom_out[158] + v_in_1[158] + e2_ext[158]};
//assign v_1[159] = {16'd0, decom_out[159] + v_in_1[159] + e2_ext[159]};
//assign v_1[160] = {16'd0, decom_out[160] + v_in_1[160] + e2_ext[160]};
//assign v_1[161] = {16'd0, decom_out[161] + v_in_1[161] + e2_ext[161]};
//assign v_1[162] = {16'd0, decom_out[162] + v_in_1[162] + e2_ext[162]};
//assign v_1[163] = {16'd0, decom_out[163] + v_in_1[163] + e2_ext[163]};
//assign v_1[164] = {16'd0, decom_out[164] + v_in_1[164] + e2_ext[164]};
//assign v_1[165] = {16'd0, decom_out[165] + v_in_1[165] + e2_ext[165]};
//assign v_1[166] = {16'd0, decom_out[166] + v_in_1[166] + e2_ext[166]};
//assign v_1[167] = {16'd0, decom_out[167] + v_in_1[167] + e2_ext[167]};
//assign v_1[168] = {16'd0, decom_out[168] + v_in_1[168] + e2_ext[168]};
//assign v_1[169] = {16'd0, decom_out[169] + v_in_1[169] + e2_ext[169]};
//assign v_1[170] = {16'd0, decom_out[170] + v_in_1[170] + e2_ext[170]};
//assign v_1[171] = {16'd0, decom_out[171] + v_in_1[171] + e2_ext[171]};
//assign v_1[172] = {16'd0, decom_out[172] + v_in_1[172] + e2_ext[172]};
//assign v_1[173] = {16'd0, decom_out[173] + v_in_1[173] + e2_ext[173]};
//assign v_1[174] = {16'd0, decom_out[174] + v_in_1[174] + e2_ext[174]};
//assign v_1[175] = {16'd0, decom_out[175] + v_in_1[175] + e2_ext[175]};
//assign v_1[176] = {16'd0, decom_out[176] + v_in_1[176] + e2_ext[176]};
//assign v_1[177] = {16'd0, decom_out[177] + v_in_1[177] + e2_ext[177]};
//assign v_1[178] = {16'd0, decom_out[178] + v_in_1[178] + e2_ext[178]};
//assign v_1[179] = {16'd0, decom_out[179] + v_in_1[179] + e2_ext[179]};
//assign v_1[180] = {16'd0, decom_out[180] + v_in_1[180] + e2_ext[180]};
//assign v_1[181] = {16'd0, decom_out[181] + v_in_1[181] + e2_ext[181]};
//assign v_1[182] = {16'd0, decom_out[182] + v_in_1[182] + e2_ext[182]};
//assign v_1[183] = {16'd0, decom_out[183] + v_in_1[183] + e2_ext[183]};
//assign v_1[184] = {16'd0, decom_out[184] + v_in_1[184] + e2_ext[184]};
//assign v_1[185] = {16'd0, decom_out[185] + v_in_1[185] + e2_ext[185]};
//assign v_1[186] = {16'd0, decom_out[186] + v_in_1[186] + e2_ext[186]};
//assign v_1[187] = {16'd0, decom_out[187] + v_in_1[187] + e2_ext[187]};
//assign v_1[188] = {16'd0, decom_out[188] + v_in_1[188] + e2_ext[188]};
//assign v_1[189] = {16'd0, decom_out[189] + v_in_1[189] + e2_ext[189]};
//assign v_1[190] = {16'd0, decom_out[190] + v_in_1[190] + e2_ext[190]};
//assign v_1[191] = {16'd0, decom_out[191] + v_in_1[191] + e2_ext[191]};
//assign v_1[192] = {16'd0, decom_out[192] + v_in_1[192] + e2_ext[192]};
//assign v_1[193] = {16'd0, decom_out[193] + v_in_1[193] + e2_ext[193]};
//assign v_1[194] = {16'd0, decom_out[194] + v_in_1[194] + e2_ext[194]};
//assign v_1[195] = {16'd0, decom_out[195] + v_in_1[195] + e2_ext[195]};
//assign v_1[196] = {16'd0, decom_out[196] + v_in_1[196] + e2_ext[196]};
//assign v_1[197] = {16'd0, decom_out[197] + v_in_1[197] + e2_ext[197]};
//assign v_1[198] = {16'd0, decom_out[198] + v_in_1[198] + e2_ext[198]};
//assign v_1[199] = {16'd0, decom_out[199] + v_in_1[199] + e2_ext[199]};
//assign v_1[200] = {16'd0, decom_out[200] + v_in_1[200] + e2_ext[200]};
//assign v_1[201] = {16'd0, decom_out[201] + v_in_1[201] + e2_ext[201]};
//assign v_1[202] = {16'd0, decom_out[202] + v_in_1[202] + e2_ext[202]};
//assign v_1[203] = {16'd0, decom_out[203] + v_in_1[203] + e2_ext[203]};
//assign v_1[204] = {16'd0, decom_out[204] + v_in_1[204] + e2_ext[204]};
//assign v_1[205] = {16'd0, decom_out[205] + v_in_1[205] + e2_ext[205]};
//assign v_1[206] = {16'd0, decom_out[206] + v_in_1[206] + e2_ext[206]};
//assign v_1[207] = {16'd0, decom_out[207] + v_in_1[207] + e2_ext[207]};
//assign v_1[208] = {16'd0, decom_out[208] + v_in_1[208] + e2_ext[208]};
//assign v_1[209] = {16'd0, decom_out[209] + v_in_1[209] + e2_ext[209]};
//assign v_1[210] = {16'd0, decom_out[210] + v_in_1[210] + e2_ext[210]};
//assign v_1[211] = {16'd0, decom_out[211] + v_in_1[211] + e2_ext[211]};
//assign v_1[212] = {16'd0, decom_out[212] + v_in_1[212] + e2_ext[212]};
//assign v_1[213] = {16'd0, decom_out[213] + v_in_1[213] + e2_ext[213]};
//assign v_1[214] = {16'd0, decom_out[214] + v_in_1[214] + e2_ext[214]};
//assign v_1[215] = {16'd0, decom_out[215] + v_in_1[215] + e2_ext[215]};
//assign v_1[216] = {16'd0, decom_out[216] + v_in_1[216] + e2_ext[216]};
//assign v_1[217] = {16'd0, decom_out[217] + v_in_1[217] + e2_ext[217]};
//assign v_1[218] = {16'd0, decom_out[218] + v_in_1[218] + e2_ext[218]};
//assign v_1[219] = {16'd0, decom_out[219] + v_in_1[219] + e2_ext[219]};
//assign v_1[220] = {16'd0, decom_out[220] + v_in_1[220] + e2_ext[220]};
//assign v_1[221] = {16'd0, decom_out[221] + v_in_1[221] + e2_ext[221]};
//assign v_1[222] = {16'd0, decom_out[222] + v_in_1[222] + e2_ext[222]};
//assign v_1[223] = {16'd0, decom_out[223] + v_in_1[223] + e2_ext[223]};
//assign v_1[224] = {16'd0, decom_out[224] + v_in_1[224] + e2_ext[224]};
//assign v_1[225] = {16'd0, decom_out[225] + v_in_1[225] + e2_ext[225]};
//assign v_1[226] = {16'd0, decom_out[226] + v_in_1[226] + e2_ext[226]};
//assign v_1[227] = {16'd0, decom_out[227] + v_in_1[227] + e2_ext[227]};
//assign v_1[228] = {16'd0, decom_out[228] + v_in_1[228] + e2_ext[228]};
//assign v_1[229] = {16'd0, decom_out[229] + v_in_1[229] + e2_ext[229]};
//assign v_1[230] = {16'd0, decom_out[230] + v_in_1[230] + e2_ext[230]};
//assign v_1[231] = {16'd0, decom_out[231] + v_in_1[231] + e2_ext[231]};
//assign v_1[232] = {16'd0, decom_out[232] + v_in_1[232] + e2_ext[232]};
//assign v_1[233] = {16'd0, decom_out[233] + v_in_1[233] + e2_ext[233]};
//assign v_1[234] = {16'd0, decom_out[234] + v_in_1[234] + e2_ext[234]};
//assign v_1[235] = {16'd0, decom_out[235] + v_in_1[235] + e2_ext[235]};
//assign v_1[236] = {16'd0, decom_out[236] + v_in_1[236] + e2_ext[236]};
//assign v_1[237] = {16'd0, decom_out[237] + v_in_1[237] + e2_ext[237]};
//assign v_1[238] = {16'd0, decom_out[238] + v_in_1[238] + e2_ext[238]};
//assign v_1[239] = {16'd0, decom_out[239] + v_in_1[239] + e2_ext[239]};
//assign v_1[240] = {16'd0, decom_out[240] + v_in_1[240] + e2_ext[240]};
//assign v_1[241] = {16'd0, decom_out[241] + v_in_1[241] + e2_ext[241]};
//assign v_1[242] = {16'd0, decom_out[242] + v_in_1[242] + e2_ext[242]};
//assign v_1[243] = {16'd0, decom_out[243] + v_in_1[243] + e2_ext[243]};
//assign v_1[244] = {16'd0, decom_out[244] + v_in_1[244] + e2_ext[244]};
//assign v_1[245] = {16'd0, decom_out[245] + v_in_1[245] + e2_ext[245]};
//assign v_1[246] = {16'd0, decom_out[246] + v_in_1[246] + e2_ext[246]};
//assign v_1[247] = {16'd0, decom_out[247] + v_in_1[247] + e2_ext[247]};
//assign v_1[248] = {16'd0, decom_out[248] + v_in_1[248] + e2_ext[248]};
//assign v_1[249] = {16'd0, decom_out[249] + v_in_1[249] + e2_ext[249]};
//assign v_1[250] = {16'd0, decom_out[250] + v_in_1[250] + e2_ext[250]};
//assign v_1[251] = {16'd0, decom_out[251] + v_in_1[251] + e2_ext[251]};
//assign v_1[252] = {16'd0, decom_out[252] + v_in_1[252] + e2_ext[252]};
//assign v_1[253] = {16'd0, decom_out[253] + v_in_1[253] + e2_ext[253]};
//assign v_1[254] = {16'd0, decom_out[254] + v_in_1[254] + e2_ext[254]};
//assign v_1[255] = {16'd0, decom_out[255] + v_in_1[255] + e2_ext[255]};

//assign v_2[0] = {16'd0, decom_out[0] + v_in_2[0] + e2_ext[0]};
//assign v_2[1] = {16'd0, decom_out[1] + v_in_2[1] + e2_ext[1]};
//assign v_2[2] = {16'd0, decom_out[2] + v_in_2[2] + e2_ext[2]};
//assign v_2[3] = {16'd0, decom_out[3] + v_in_2[3] + e2_ext[3]};
//assign v_2[4] = {16'd0, decom_out[4] + v_in_2[4] + e2_ext[4]};
//assign v_2[5] = {16'd0, decom_out[5] + v_in_2[5] + e2_ext[5]};
//assign v_2[6] = {16'd0, decom_out[6] + v_in_2[6] + e2_ext[6]};
//assign v_2[7] = {16'd0, decom_out[7] + v_in_2[7] + e2_ext[7]};
//assign v_2[8] = {16'd0, decom_out[8] + v_in_2[8] + e2_ext[8]};
//assign v_2[9] = {16'd0, decom_out[9] + v_in_2[9] + e2_ext[9]};
//assign v_2[10] = {16'd0, decom_out[10] + v_in_2[10] + e2_ext[10]};
//assign v_2[11] = {16'd0, decom_out[11] + v_in_2[11] + e2_ext[11]};
//assign v_2[12] = {16'd0, decom_out[12] + v_in_2[12] + e2_ext[12]};
//assign v_2[13] = {16'd0, decom_out[13] + v_in_2[13] + e2_ext[13]};
//assign v_2[14] = {16'd0, decom_out[14] + v_in_2[14] + e2_ext[14]};
//assign v_2[15] = {16'd0, decom_out[15] + v_in_2[15] + e2_ext[15]};
//assign v_2[16] = {16'd0, decom_out[16] + v_in_2[16] + e2_ext[16]};
//assign v_2[17] = {16'd0, decom_out[17] + v_in_2[17] + e2_ext[17]};
//assign v_2[18] = {16'd0, decom_out[18] + v_in_2[18] + e2_ext[18]};
//assign v_2[19] = {16'd0, decom_out[19] + v_in_2[19] + e2_ext[19]};
//assign v_2[20] = {16'd0, decom_out[20] + v_in_2[20] + e2_ext[20]};
//assign v_2[21] = {16'd0, decom_out[21] + v_in_2[21] + e2_ext[21]};
//assign v_2[22] = {16'd0, decom_out[22] + v_in_2[22] + e2_ext[22]};
//assign v_2[23] = {16'd0, decom_out[23] + v_in_2[23] + e2_ext[23]};
//assign v_2[24] = {16'd0, decom_out[24] + v_in_2[24] + e2_ext[24]};
//assign v_2[25] = {16'd0, decom_out[25] + v_in_2[25] + e2_ext[25]};
//assign v_2[26] = {16'd0, decom_out[26] + v_in_2[26] + e2_ext[26]};
//assign v_2[27] = {16'd0, decom_out[27] + v_in_2[27] + e2_ext[27]};
//assign v_2[28] = {16'd0, decom_out[28] + v_in_2[28] + e2_ext[28]};
//assign v_2[29] = {16'd0, decom_out[29] + v_in_2[29] + e2_ext[29]};
//assign v_2[30] = {16'd0, decom_out[30] + v_in_2[30] + e2_ext[30]};
//assign v_2[31] = {16'd0, decom_out[31] + v_in_2[31] + e2_ext[31]};
//assign v_2[32] = {16'd0, decom_out[32] + v_in_2[32] + e2_ext[32]};
//assign v_2[33] = {16'd0, decom_out[33] + v_in_2[33] + e2_ext[33]};
//assign v_2[34] = {16'd0, decom_out[34] + v_in_2[34] + e2_ext[34]};
//assign v_2[35] = {16'd0, decom_out[35] + v_in_2[35] + e2_ext[35]};
//assign v_2[36] = {16'd0, decom_out[36] + v_in_2[36] + e2_ext[36]};
//assign v_2[37] = {16'd0, decom_out[37] + v_in_2[37] + e2_ext[37]};
//assign v_2[38] = {16'd0, decom_out[38] + v_in_2[38] + e2_ext[38]};
//assign v_2[39] = {16'd0, decom_out[39] + v_in_2[39] + e2_ext[39]};
//assign v_2[40] = {16'd0, decom_out[40] + v_in_2[40] + e2_ext[40]};
//assign v_2[41] = {16'd0, decom_out[41] + v_in_2[41] + e2_ext[41]};
//assign v_2[42] = {16'd0, decom_out[42] + v_in_2[42] + e2_ext[42]};
//assign v_2[43] = {16'd0, decom_out[43] + v_in_2[43] + e2_ext[43]};
//assign v_2[44] = {16'd0, decom_out[44] + v_in_2[44] + e2_ext[44]};
//assign v_2[45] = {16'd0, decom_out[45] + v_in_2[45] + e2_ext[45]};
//assign v_2[46] = {16'd0, decom_out[46] + v_in_2[46] + e2_ext[46]};
//assign v_2[47] = {16'd0, decom_out[47] + v_in_2[47] + e2_ext[47]};
//assign v_2[48] = {16'd0, decom_out[48] + v_in_2[48] + e2_ext[48]};
//assign v_2[49] = {16'd0, decom_out[49] + v_in_2[49] + e2_ext[49]};
//assign v_2[50] = {16'd0, decom_out[50] + v_in_2[50] + e2_ext[50]};
//assign v_2[51] = {16'd0, decom_out[51] + v_in_2[51] + e2_ext[51]};
//assign v_2[52] = {16'd0, decom_out[52] + v_in_2[52] + e2_ext[52]};
//assign v_2[53] = {16'd0, decom_out[53] + v_in_2[53] + e2_ext[53]};
//assign v_2[54] = {16'd0, decom_out[54] + v_in_2[54] + e2_ext[54]};
//assign v_2[55] = {16'd0, decom_out[55] + v_in_2[55] + e2_ext[55]};
//assign v_2[56] = {16'd0, decom_out[56] + v_in_2[56] + e2_ext[56]};
//assign v_2[57] = {16'd0, decom_out[57] + v_in_2[57] + e2_ext[57]};
//assign v_2[58] = {16'd0, decom_out[58] + v_in_2[58] + e2_ext[58]};
//assign v_2[59] = {16'd0, decom_out[59] + v_in_2[59] + e2_ext[59]};
//assign v_2[60] = {16'd0, decom_out[60] + v_in_2[60] + e2_ext[60]};
//assign v_2[61] = {16'd0, decom_out[61] + v_in_2[61] + e2_ext[61]};
//assign v_2[62] = {16'd0, decom_out[62] + v_in_2[62] + e2_ext[62]};
//assign v_2[63] = {16'd0, decom_out[63] + v_in_2[63] + e2_ext[63]};
//assign v_2[64] = {16'd0, decom_out[64] + v_in_2[64] + e2_ext[64]};
//assign v_2[65] = {16'd0, decom_out[65] + v_in_2[65] + e2_ext[65]};
//assign v_2[66] = {16'd0, decom_out[66] + v_in_2[66] + e2_ext[66]};
//assign v_2[67] = {16'd0, decom_out[67] + v_in_2[67] + e2_ext[67]};
//assign v_2[68] = {16'd0, decom_out[68] + v_in_2[68] + e2_ext[68]};
//assign v_2[69] = {16'd0, decom_out[69] + v_in_2[69] + e2_ext[69]};
//assign v_2[70] = {16'd0, decom_out[70] + v_in_2[70] + e2_ext[70]};
//assign v_2[71] = {16'd0, decom_out[71] + v_in_2[71] + e2_ext[71]};
//assign v_2[72] = {16'd0, decom_out[72] + v_in_2[72] + e2_ext[72]};
//assign v_2[73] = {16'd0, decom_out[73] + v_in_2[73] + e2_ext[73]};
//assign v_2[74] = {16'd0, decom_out[74] + v_in_2[74] + e2_ext[74]};
//assign v_2[75] = {16'd0, decom_out[75] + v_in_2[75] + e2_ext[75]};
//assign v_2[76] = {16'd0, decom_out[76] + v_in_2[76] + e2_ext[76]};
//assign v_2[77] = {16'd0, decom_out[77] + v_in_2[77] + e2_ext[77]};
//assign v_2[78] = {16'd0, decom_out[78] + v_in_2[78] + e2_ext[78]};
//assign v_2[79] = {16'd0, decom_out[79] + v_in_2[79] + e2_ext[79]};
//assign v_2[80] = {16'd0, decom_out[80] + v_in_2[80] + e2_ext[80]};
//assign v_2[81] = {16'd0, decom_out[81] + v_in_2[81] + e2_ext[81]};
//assign v_2[82] = {16'd0, decom_out[82] + v_in_2[82] + e2_ext[82]};
//assign v_2[83] = {16'd0, decom_out[83] + v_in_2[83] + e2_ext[83]};
//assign v_2[84] = {16'd0, decom_out[84] + v_in_2[84] + e2_ext[84]};
//assign v_2[85] = {16'd0, decom_out[85] + v_in_2[85] + e2_ext[85]};
//assign v_2[86] = {16'd0, decom_out[86] + v_in_2[86] + e2_ext[86]};
//assign v_2[87] = {16'd0, decom_out[87] + v_in_2[87] + e2_ext[87]};
//assign v_2[88] = {16'd0, decom_out[88] + v_in_2[88] + e2_ext[88]};
//assign v_2[89] = {16'd0, decom_out[89] + v_in_2[89] + e2_ext[89]};
//assign v_2[90] = {16'd0, decom_out[90] + v_in_2[90] + e2_ext[90]};
//assign v_2[91] = {16'd0, decom_out[91] + v_in_2[91] + e2_ext[91]};
//assign v_2[92] = {16'd0, decom_out[92] + v_in_2[92] + e2_ext[92]};
//assign v_2[93] = {16'd0, decom_out[93] + v_in_2[93] + e2_ext[93]};
//assign v_2[94] = {16'd0, decom_out[94] + v_in_2[94] + e2_ext[94]};
//assign v_2[95] = {16'd0, decom_out[95] + v_in_2[95] + e2_ext[95]};
//assign v_2[96] = {16'd0, decom_out[96] + v_in_2[96] + e2_ext[96]};
//assign v_2[97] = {16'd0, decom_out[97] + v_in_2[97] + e2_ext[97]};
//assign v_2[98] = {16'd0, decom_out[98] + v_in_2[98] + e2_ext[98]};
//assign v_2[99] = {16'd0, decom_out[99] + v_in_2[99] + e2_ext[99]};
//assign v_2[100] = {16'd0, decom_out[100] + v_in_2[100] + e2_ext[100]};
//assign v_2[101] = {16'd0, decom_out[101] + v_in_2[101] + e2_ext[101]};
//assign v_2[102] = {16'd0, decom_out[102] + v_in_2[102] + e2_ext[102]};
//assign v_2[103] = {16'd0, decom_out[103] + v_in_2[103] + e2_ext[103]};
//assign v_2[104] = {16'd0, decom_out[104] + v_in_2[104] + e2_ext[104]};
//assign v_2[105] = {16'd0, decom_out[105] + v_in_2[105] + e2_ext[105]};
//assign v_2[106] = {16'd0, decom_out[106] + v_in_2[106] + e2_ext[106]};
//assign v_2[107] = {16'd0, decom_out[107] + v_in_2[107] + e2_ext[107]};
//assign v_2[108] = {16'd0, decom_out[108] + v_in_2[108] + e2_ext[108]};
//assign v_2[109] = {16'd0, decom_out[109] + v_in_2[109] + e2_ext[109]};
//assign v_2[110] = {16'd0, decom_out[110] + v_in_2[110] + e2_ext[110]};
//assign v_2[111] = {16'd0, decom_out[111] + v_in_2[111] + e2_ext[111]};
//assign v_2[112] = {16'd0, decom_out[112] + v_in_2[112] + e2_ext[112]};
//assign v_2[113] = {16'd0, decom_out[113] + v_in_2[113] + e2_ext[113]};
//assign v_2[114] = {16'd0, decom_out[114] + v_in_2[114] + e2_ext[114]};
//assign v_2[115] = {16'd0, decom_out[115] + v_in_2[115] + e2_ext[115]};
//assign v_2[116] = {16'd0, decom_out[116] + v_in_2[116] + e2_ext[116]};
//assign v_2[117] = {16'd0, decom_out[117] + v_in_2[117] + e2_ext[117]};
//assign v_2[118] = {16'd0, decom_out[118] + v_in_2[118] + e2_ext[118]};
//assign v_2[119] = {16'd0, decom_out[119] + v_in_2[119] + e2_ext[119]};
//assign v_2[120] = {16'd0, decom_out[120] + v_in_2[120] + e2_ext[120]};
//assign v_2[121] = {16'd0, decom_out[121] + v_in_2[121] + e2_ext[121]};
//assign v_2[122] = {16'd0, decom_out[122] + v_in_2[122] + e2_ext[122]};
//assign v_2[123] = {16'd0, decom_out[123] + v_in_2[123] + e2_ext[123]};
//assign v_2[124] = {16'd0, decom_out[124] + v_in_2[124] + e2_ext[124]};
//assign v_2[125] = {16'd0, decom_out[125] + v_in_2[125] + e2_ext[125]};
//assign v_2[126] = {16'd0, decom_out[126] + v_in_2[126] + e2_ext[126]};
//assign v_2[127] = {16'd0, decom_out[127] + v_in_2[127] + e2_ext[127]};
//assign v_2[128] = {16'd0, decom_out[128] + v_in_2[128] + e2_ext[128]};
//assign v_2[129] = {16'd0, decom_out[129] + v_in_2[129] + e2_ext[129]};
//assign v_2[130] = {16'd0, decom_out[130] + v_in_2[130] + e2_ext[130]};
//assign v_2[131] = {16'd0, decom_out[131] + v_in_2[131] + e2_ext[131]};
//assign v_2[132] = {16'd0, decom_out[132] + v_in_2[132] + e2_ext[132]};
//assign v_2[133] = {16'd0, decom_out[133] + v_in_2[133] + e2_ext[133]};
//assign v_2[134] = {16'd0, decom_out[134] + v_in_2[134] + e2_ext[134]};
//assign v_2[135] = {16'd0, decom_out[135] + v_in_2[135] + e2_ext[135]};
//assign v_2[136] = {16'd0, decom_out[136] + v_in_2[136] + e2_ext[136]};
//assign v_2[137] = {16'd0, decom_out[137] + v_in_2[137] + e2_ext[137]};
//assign v_2[138] = {16'd0, decom_out[138] + v_in_2[138] + e2_ext[138]};
//assign v_2[139] = {16'd0, decom_out[139] + v_in_2[139] + e2_ext[139]};
//assign v_2[140] = {16'd0, decom_out[140] + v_in_2[140] + e2_ext[140]};
//assign v_2[141] = {16'd0, decom_out[141] + v_in_2[141] + e2_ext[141]};
//assign v_2[142] = {16'd0, decom_out[142] + v_in_2[142] + e2_ext[142]};
//assign v_2[143] = {16'd0, decom_out[143] + v_in_2[143] + e2_ext[143]};
//assign v_2[144] = {16'd0, decom_out[144] + v_in_2[144] + e2_ext[144]};
//assign v_2[145] = {16'd0, decom_out[145] + v_in_2[145] + e2_ext[145]};
//assign v_2[146] = {16'd0, decom_out[146] + v_in_2[146] + e2_ext[146]};
//assign v_2[147] = {16'd0, decom_out[147] + v_in_2[147] + e2_ext[147]};
//assign v_2[148] = {16'd0, decom_out[148] + v_in_2[148] + e2_ext[148]};
//assign v_2[149] = {16'd0, decom_out[149] + v_in_2[149] + e2_ext[149]};
//assign v_2[150] = {16'd0, decom_out[150] + v_in_2[150] + e2_ext[150]};
//assign v_2[151] = {16'd0, decom_out[151] + v_in_2[151] + e2_ext[151]};
//assign v_2[152] = {16'd0, decom_out[152] + v_in_2[152] + e2_ext[152]};
//assign v_2[153] = {16'd0, decom_out[153] + v_in_2[153] + e2_ext[153]};
//assign v_2[154] = {16'd0, decom_out[154] + v_in_2[154] + e2_ext[154]};
//assign v_2[155] = {16'd0, decom_out[155] + v_in_2[155] + e2_ext[155]};
//assign v_2[156] = {16'd0, decom_out[156] + v_in_2[156] + e2_ext[156]};
//assign v_2[157] = {16'd0, decom_out[157] + v_in_2[157] + e2_ext[157]};
//assign v_2[158] = {16'd0, decom_out[158] + v_in_2[158] + e2_ext[158]};
//assign v_2[159] = {16'd0, decom_out[159] + v_in_2[159] + e2_ext[159]};
//assign v_2[160] = {16'd0, decom_out[160] + v_in_2[160] + e2_ext[160]};
//assign v_2[161] = {16'd0, decom_out[161] + v_in_2[161] + e2_ext[161]};
//assign v_2[162] = {16'd0, decom_out[162] + v_in_2[162] + e2_ext[162]};
//assign v_2[163] = {16'd0, decom_out[163] + v_in_2[163] + e2_ext[163]};
//assign v_2[164] = {16'd0, decom_out[164] + v_in_2[164] + e2_ext[164]};
//assign v_2[165] = {16'd0, decom_out[165] + v_in_2[165] + e2_ext[165]};
//assign v_2[166] = {16'd0, decom_out[166] + v_in_2[166] + e2_ext[166]};
//assign v_2[167] = {16'd0, decom_out[167] + v_in_2[167] + e2_ext[167]};
//assign v_2[168] = {16'd0, decom_out[168] + v_in_2[168] + e2_ext[168]};
//assign v_2[169] = {16'd0, decom_out[169] + v_in_2[169] + e2_ext[169]};
//assign v_2[170] = {16'd0, decom_out[170] + v_in_2[170] + e2_ext[170]};
//assign v_2[171] = {16'd0, decom_out[171] + v_in_2[171] + e2_ext[171]};
//assign v_2[172] = {16'd0, decom_out[172] + v_in_2[172] + e2_ext[172]};
//assign v_2[173] = {16'd0, decom_out[173] + v_in_2[173] + e2_ext[173]};
//assign v_2[174] = {16'd0, decom_out[174] + v_in_2[174] + e2_ext[174]};
//assign v_2[175] = {16'd0, decom_out[175] + v_in_2[175] + e2_ext[175]};
//assign v_2[176] = {16'd0, decom_out[176] + v_in_2[176] + e2_ext[176]};
//assign v_2[177] = {16'd0, decom_out[177] + v_in_2[177] + e2_ext[177]};
//assign v_2[178] = {16'd0, decom_out[178] + v_in_2[178] + e2_ext[178]};
//assign v_2[179] = {16'd0, decom_out[179] + v_in_2[179] + e2_ext[179]};
//assign v_2[180] = {16'd0, decom_out[180] + v_in_2[180] + e2_ext[180]};
//assign v_2[181] = {16'd0, decom_out[181] + v_in_2[181] + e2_ext[181]};
//assign v_2[182] = {16'd0, decom_out[182] + v_in_2[182] + e2_ext[182]};
//assign v_2[183] = {16'd0, decom_out[183] + v_in_2[183] + e2_ext[183]};
//assign v_2[184] = {16'd0, decom_out[184] + v_in_2[184] + e2_ext[184]};
//assign v_2[185] = {16'd0, decom_out[185] + v_in_2[185] + e2_ext[185]};
//assign v_2[186] = {16'd0, decom_out[186] + v_in_2[186] + e2_ext[186]};
//assign v_2[187] = {16'd0, decom_out[187] + v_in_2[187] + e2_ext[187]};
//assign v_2[188] = {16'd0, decom_out[188] + v_in_2[188] + e2_ext[188]};
//assign v_2[189] = {16'd0, decom_out[189] + v_in_2[189] + e2_ext[189]};
//assign v_2[190] = {16'd0, decom_out[190] + v_in_2[190] + e2_ext[190]};
//assign v_2[191] = {16'd0, decom_out[191] + v_in_2[191] + e2_ext[191]};
//assign v_2[192] = {16'd0, decom_out[192] + v_in_2[192] + e2_ext[192]};
//assign v_2[193] = {16'd0, decom_out[193] + v_in_2[193] + e2_ext[193]};
//assign v_2[194] = {16'd0, decom_out[194] + v_in_2[194] + e2_ext[194]};
//assign v_2[195] = {16'd0, decom_out[195] + v_in_2[195] + e2_ext[195]};
//assign v_2[196] = {16'd0, decom_out[196] + v_in_2[196] + e2_ext[196]};
//assign v_2[197] = {16'd0, decom_out[197] + v_in_2[197] + e2_ext[197]};
//assign v_2[198] = {16'd0, decom_out[198] + v_in_2[198] + e2_ext[198]};
//assign v_2[199] = {16'd0, decom_out[199] + v_in_2[199] + e2_ext[199]};
//assign v_2[200] = {16'd0, decom_out[200] + v_in_2[200] + e2_ext[200]};
//assign v_2[201] = {16'd0, decom_out[201] + v_in_2[201] + e2_ext[201]};
//assign v_2[202] = {16'd0, decom_out[202] + v_in_2[202] + e2_ext[202]};
//assign v_2[203] = {16'd0, decom_out[203] + v_in_2[203] + e2_ext[203]};
//assign v_2[204] = {16'd0, decom_out[204] + v_in_2[204] + e2_ext[204]};
//assign v_2[205] = {16'd0, decom_out[205] + v_in_2[205] + e2_ext[205]};
//assign v_2[206] = {16'd0, decom_out[206] + v_in_2[206] + e2_ext[206]};
//assign v_2[207] = {16'd0, decom_out[207] + v_in_2[207] + e2_ext[207]};
//assign v_2[208] = {16'd0, decom_out[208] + v_in_2[208] + e2_ext[208]};
//assign v_2[209] = {16'd0, decom_out[209] + v_in_2[209] + e2_ext[209]};
//assign v_2[210] = {16'd0, decom_out[210] + v_in_2[210] + e2_ext[210]};
//assign v_2[211] = {16'd0, decom_out[211] + v_in_2[211] + e2_ext[211]};
//assign v_2[212] = {16'd0, decom_out[212] + v_in_2[212] + e2_ext[212]};
//assign v_2[213] = {16'd0, decom_out[213] + v_in_2[213] + e2_ext[213]};
//assign v_2[214] = {16'd0, decom_out[214] + v_in_2[214] + e2_ext[214]};
//assign v_2[215] = {16'd0, decom_out[215] + v_in_2[215] + e2_ext[215]};
//assign v_2[216] = {16'd0, decom_out[216] + v_in_2[216] + e2_ext[216]};
//assign v_2[217] = {16'd0, decom_out[217] + v_in_2[217] + e2_ext[217]};
//assign v_2[218] = {16'd0, decom_out[218] + v_in_2[218] + e2_ext[218]};
//assign v_2[219] = {16'd0, decom_out[219] + v_in_2[219] + e2_ext[219]};
//assign v_2[220] = {16'd0, decom_out[220] + v_in_2[220] + e2_ext[220]};
//assign v_2[221] = {16'd0, decom_out[221] + v_in_2[221] + e2_ext[221]};
//assign v_2[222] = {16'd0, decom_out[222] + v_in_2[222] + e2_ext[222]};
//assign v_2[223] = {16'd0, decom_out[223] + v_in_2[223] + e2_ext[223]};
//assign v_2[224] = {16'd0, decom_out[224] + v_in_2[224] + e2_ext[224]};
//assign v_2[225] = {16'd0, decom_out[225] + v_in_2[225] + e2_ext[225]};
//assign v_2[226] = {16'd0, decom_out[226] + v_in_2[226] + e2_ext[226]};
//assign v_2[227] = {16'd0, decom_out[227] + v_in_2[227] + e2_ext[227]};
//assign v_2[228] = {16'd0, decom_out[228] + v_in_2[228] + e2_ext[228]};
//assign v_2[229] = {16'd0, decom_out[229] + v_in_2[229] + e2_ext[229]};
//assign v_2[230] = {16'd0, decom_out[230] + v_in_2[230] + e2_ext[230]};
//assign v_2[231] = {16'd0, decom_out[231] + v_in_2[231] + e2_ext[231]};
//assign v_2[232] = {16'd0, decom_out[232] + v_in_2[232] + e2_ext[232]};
//assign v_2[233] = {16'd0, decom_out[233] + v_in_2[233] + e2_ext[233]};
//assign v_2[234] = {16'd0, decom_out[234] + v_in_2[234] + e2_ext[234]};
//assign v_2[235] = {16'd0, decom_out[235] + v_in_2[235] + e2_ext[235]};
//assign v_2[236] = {16'd0, decom_out[236] + v_in_2[236] + e2_ext[236]};
//assign v_2[237] = {16'd0, decom_out[237] + v_in_2[237] + e2_ext[237]};
//assign v_2[238] = {16'd0, decom_out[238] + v_in_2[238] + e2_ext[238]};
//assign v_2[239] = {16'd0, decom_out[239] + v_in_2[239] + e2_ext[239]};
//assign v_2[240] = {16'd0, decom_out[240] + v_in_2[240] + e2_ext[240]};
//assign v_2[241] = {16'd0, decom_out[241] + v_in_2[241] + e2_ext[241]};
//assign v_2[242] = {16'd0, decom_out[242] + v_in_2[242] + e2_ext[242]};
//assign v_2[243] = {16'd0, decom_out[243] + v_in_2[243] + e2_ext[243]};
//assign v_2[244] = {16'd0, decom_out[244] + v_in_2[244] + e2_ext[244]};
//assign v_2[245] = {16'd0, decom_out[245] + v_in_2[245] + e2_ext[245]};
//assign v_2[246] = {16'd0, decom_out[246] + v_in_2[246] + e2_ext[246]};
//assign v_2[247] = {16'd0, decom_out[247] + v_in_2[247] + e2_ext[247]};
//assign v_2[248] = {16'd0, decom_out[248] + v_in_2[248] + e2_ext[248]};
//assign v_2[249] = {16'd0, decom_out[249] + v_in_2[249] + e2_ext[249]};
//assign v_2[250] = {16'd0, decom_out[250] + v_in_2[250] + e2_ext[250]};
//assign v_2[251] = {16'd0, decom_out[251] + v_in_2[251] + e2_ext[251]};
//assign v_2[252] = {16'd0, decom_out[252] + v_in_2[252] + e2_ext[252]};
//assign v_2[253] = {16'd0, decom_out[253] + v_in_2[253] + e2_ext[253]};
//assign v_2[254] = {16'd0, decom_out[254] + v_in_2[254] + e2_ext[254]};
//assign v_2[255] = {16'd0, decom_out[255] + v_in_2[255] + e2_ext[255]};

//assign v_3[0] = {16'd0, decom_out[0] + v_in_3[0] + e2_ext[0]};
//assign v_3[1] = {16'd0, decom_out[1] + v_in_3[1] + e2_ext[1]};
//assign v_3[2] = {16'd0, decom_out[2] + v_in_3[2] + e2_ext[2]};
//assign v_3[3] = {16'd0, decom_out[3] + v_in_3[3] + e2_ext[3]};
//assign v_3[4] = {16'd0, decom_out[4] + v_in_3[4] + e2_ext[4]};
//assign v_3[5] = {16'd0, decom_out[5] + v_in_3[5] + e2_ext[5]};
//assign v_3[6] = {16'd0, decom_out[6] + v_in_3[6] + e2_ext[6]};
//assign v_3[7] = {16'd0, decom_out[7] + v_in_3[7] + e2_ext[7]};
//assign v_3[8] = {16'd0, decom_out[8] + v_in_3[8] + e2_ext[8]};
//assign v_3[9] = {16'd0, decom_out[9] + v_in_3[9] + e2_ext[9]};
//assign v_3[10] = {16'd0, decom_out[10] + v_in_3[10] + e2_ext[10]};
//assign v_3[11] = {16'd0, decom_out[11] + v_in_3[11] + e2_ext[11]};
//assign v_3[12] = {16'd0, decom_out[12] + v_in_3[12] + e2_ext[12]};
//assign v_3[13] = {16'd0, decom_out[13] + v_in_3[13] + e2_ext[13]};
//assign v_3[14] = {16'd0, decom_out[14] + v_in_3[14] + e2_ext[14]};
//assign v_3[15] = {16'd0, decom_out[15] + v_in_3[15] + e2_ext[15]};
//assign v_3[16] = {16'd0, decom_out[16] + v_in_3[16] + e2_ext[16]};
//assign v_3[17] = {16'd0, decom_out[17] + v_in_3[17] + e2_ext[17]};
//assign v_3[18] = {16'd0, decom_out[18] + v_in_3[18] + e2_ext[18]};
//assign v_3[19] = {16'd0, decom_out[19] + v_in_3[19] + e2_ext[19]};
//assign v_3[20] = {16'd0, decom_out[20] + v_in_3[20] + e2_ext[20]};
//assign v_3[21] = {16'd0, decom_out[21] + v_in_3[21] + e2_ext[21]};
//assign v_3[22] = {16'd0, decom_out[22] + v_in_3[22] + e2_ext[22]};
//assign v_3[23] = {16'd0, decom_out[23] + v_in_3[23] + e2_ext[23]};
//assign v_3[24] = {16'd0, decom_out[24] + v_in_3[24] + e2_ext[24]};
//assign v_3[25] = {16'd0, decom_out[25] + v_in_3[25] + e2_ext[25]};
//assign v_3[26] = {16'd0, decom_out[26] + v_in_3[26] + e2_ext[26]};
//assign v_3[27] = {16'd0, decom_out[27] + v_in_3[27] + e2_ext[27]};
//assign v_3[28] = {16'd0, decom_out[28] + v_in_3[28] + e2_ext[28]};
//assign v_3[29] = {16'd0, decom_out[29] + v_in_3[29] + e2_ext[29]};
//assign v_3[30] = {16'd0, decom_out[30] + v_in_3[30] + e2_ext[30]};
//assign v_3[31] = {16'd0, decom_out[31] + v_in_3[31] + e2_ext[31]};
//assign v_3[32] = {16'd0, decom_out[32] + v_in_3[32] + e2_ext[32]};
//assign v_3[33] = {16'd0, decom_out[33] + v_in_3[33] + e2_ext[33]};
//assign v_3[34] = {16'd0, decom_out[34] + v_in_3[34] + e2_ext[34]};
//assign v_3[35] = {16'd0, decom_out[35] + v_in_3[35] + e2_ext[35]};
//assign v_3[36] = {16'd0, decom_out[36] + v_in_3[36] + e2_ext[36]};
//assign v_3[37] = {16'd0, decom_out[37] + v_in_3[37] + e2_ext[37]};
//assign v_3[38] = {16'd0, decom_out[38] + v_in_3[38] + e2_ext[38]};
//assign v_3[39] = {16'd0, decom_out[39] + v_in_3[39] + e2_ext[39]};
//assign v_3[40] = {16'd0, decom_out[40] + v_in_3[40] + e2_ext[40]};
//assign v_3[41] = {16'd0, decom_out[41] + v_in_3[41] + e2_ext[41]};
//assign v_3[42] = {16'd0, decom_out[42] + v_in_3[42] + e2_ext[42]};
//assign v_3[43] = {16'd0, decom_out[43] + v_in_3[43] + e2_ext[43]};
//assign v_3[44] = {16'd0, decom_out[44] + v_in_3[44] + e2_ext[44]};
//assign v_3[45] = {16'd0, decom_out[45] + v_in_3[45] + e2_ext[45]};
//assign v_3[46] = {16'd0, decom_out[46] + v_in_3[46] + e2_ext[46]};
//assign v_3[47] = {16'd0, decom_out[47] + v_in_3[47] + e2_ext[47]};
//assign v_3[48] = {16'd0, decom_out[48] + v_in_3[48] + e2_ext[48]};
//assign v_3[49] = {16'd0, decom_out[49] + v_in_3[49] + e2_ext[49]};
//assign v_3[50] = {16'd0, decom_out[50] + v_in_3[50] + e2_ext[50]};
//assign v_3[51] = {16'd0, decom_out[51] + v_in_3[51] + e2_ext[51]};
//assign v_3[52] = {16'd0, decom_out[52] + v_in_3[52] + e2_ext[52]};
//assign v_3[53] = {16'd0, decom_out[53] + v_in_3[53] + e2_ext[53]};
//assign v_3[54] = {16'd0, decom_out[54] + v_in_3[54] + e2_ext[54]};
//assign v_3[55] = {16'd0, decom_out[55] + v_in_3[55] + e2_ext[55]};
//assign v_3[56] = {16'd0, decom_out[56] + v_in_3[56] + e2_ext[56]};
//assign v_3[57] = {16'd0, decom_out[57] + v_in_3[57] + e2_ext[57]};
//assign v_3[58] = {16'd0, decom_out[58] + v_in_3[58] + e2_ext[58]};
//assign v_3[59] = {16'd0, decom_out[59] + v_in_3[59] + e2_ext[59]};
//assign v_3[60] = {16'd0, decom_out[60] + v_in_3[60] + e2_ext[60]};
//assign v_3[61] = {16'd0, decom_out[61] + v_in_3[61] + e2_ext[61]};
//assign v_3[62] = {16'd0, decom_out[62] + v_in_3[62] + e2_ext[62]};
//assign v_3[63] = {16'd0, decom_out[63] + v_in_3[63] + e2_ext[63]};
//assign v_3[64] = {16'd0, decom_out[64] + v_in_3[64] + e2_ext[64]};
//assign v_3[65] = {16'd0, decom_out[65] + v_in_3[65] + e2_ext[65]};
//assign v_3[66] = {16'd0, decom_out[66] + v_in_3[66] + e2_ext[66]};
//assign v_3[67] = {16'd0, decom_out[67] + v_in_3[67] + e2_ext[67]};
//assign v_3[68] = {16'd0, decom_out[68] + v_in_3[68] + e2_ext[68]};
//assign v_3[69] = {16'd0, decom_out[69] + v_in_3[69] + e2_ext[69]};
//assign v_3[70] = {16'd0, decom_out[70] + v_in_3[70] + e2_ext[70]};
//assign v_3[71] = {16'd0, decom_out[71] + v_in_3[71] + e2_ext[71]};
//assign v_3[72] = {16'd0, decom_out[72] + v_in_3[72] + e2_ext[72]};
//assign v_3[73] = {16'd0, decom_out[73] + v_in_3[73] + e2_ext[73]};
//assign v_3[74] = {16'd0, decom_out[74] + v_in_3[74] + e2_ext[74]};
//assign v_3[75] = {16'd0, decom_out[75] + v_in_3[75] + e2_ext[75]};
//assign v_3[76] = {16'd0, decom_out[76] + v_in_3[76] + e2_ext[76]};
//assign v_3[77] = {16'd0, decom_out[77] + v_in_3[77] + e2_ext[77]};
//assign v_3[78] = {16'd0, decom_out[78] + v_in_3[78] + e2_ext[78]};
//assign v_3[79] = {16'd0, decom_out[79] + v_in_3[79] + e2_ext[79]};
//assign v_3[80] = {16'd0, decom_out[80] + v_in_3[80] + e2_ext[80]};
//assign v_3[81] = {16'd0, decom_out[81] + v_in_3[81] + e2_ext[81]};
//assign v_3[82] = {16'd0, decom_out[82] + v_in_3[82] + e2_ext[82]};
//assign v_3[83] = {16'd0, decom_out[83] + v_in_3[83] + e2_ext[83]};
//assign v_3[84] = {16'd0, decom_out[84] + v_in_3[84] + e2_ext[84]};
//assign v_3[85] = {16'd0, decom_out[85] + v_in_3[85] + e2_ext[85]};
//assign v_3[86] = {16'd0, decom_out[86] + v_in_3[86] + e2_ext[86]};
//assign v_3[87] = {16'd0, decom_out[87] + v_in_3[87] + e2_ext[87]};
//assign v_3[88] = {16'd0, decom_out[88] + v_in_3[88] + e2_ext[88]};
//assign v_3[89] = {16'd0, decom_out[89] + v_in_3[89] + e2_ext[89]};
//assign v_3[90] = {16'd0, decom_out[90] + v_in_3[90] + e2_ext[90]};
//assign v_3[91] = {16'd0, decom_out[91] + v_in_3[91] + e2_ext[91]};
//assign v_3[92] = {16'd0, decom_out[92] + v_in_3[92] + e2_ext[92]};
//assign v_3[93] = {16'd0, decom_out[93] + v_in_3[93] + e2_ext[93]};
//assign v_3[94] = {16'd0, decom_out[94] + v_in_3[94] + e2_ext[94]};
//assign v_3[95] = {16'd0, decom_out[95] + v_in_3[95] + e2_ext[95]};
//assign v_3[96] = {16'd0, decom_out[96] + v_in_3[96] + e2_ext[96]};
//assign v_3[97] = {16'd0, decom_out[97] + v_in_3[97] + e2_ext[97]};
//assign v_3[98] = {16'd0, decom_out[98] + v_in_3[98] + e2_ext[98]};
//assign v_3[99] = {16'd0, decom_out[99] + v_in_3[99] + e2_ext[99]};
//assign v_3[100] = {16'd0, decom_out[100] + v_in_3[100] + e2_ext[100]};
//assign v_3[101] = {16'd0, decom_out[101] + v_in_3[101] + e2_ext[101]};
//assign v_3[102] = {16'd0, decom_out[102] + v_in_3[102] + e2_ext[102]};
//assign v_3[103] = {16'd0, decom_out[103] + v_in_3[103] + e2_ext[103]};
//assign v_3[104] = {16'd0, decom_out[104] + v_in_3[104] + e2_ext[104]};
//assign v_3[105] = {16'd0, decom_out[105] + v_in_3[105] + e2_ext[105]};
//assign v_3[106] = {16'd0, decom_out[106] + v_in_3[106] + e2_ext[106]};
//assign v_3[107] = {16'd0, decom_out[107] + v_in_3[107] + e2_ext[107]};
//assign v_3[108] = {16'd0, decom_out[108] + v_in_3[108] + e2_ext[108]};
//assign v_3[109] = {16'd0, decom_out[109] + v_in_3[109] + e2_ext[109]};
//assign v_3[110] = {16'd0, decom_out[110] + v_in_3[110] + e2_ext[110]};
//assign v_3[111] = {16'd0, decom_out[111] + v_in_3[111] + e2_ext[111]};
//assign v_3[112] = {16'd0, decom_out[112] + v_in_3[112] + e2_ext[112]};
//assign v_3[113] = {16'd0, decom_out[113] + v_in_3[113] + e2_ext[113]};
//assign v_3[114] = {16'd0, decom_out[114] + v_in_3[114] + e2_ext[114]};
//assign v_3[115] = {16'd0, decom_out[115] + v_in_3[115] + e2_ext[115]};
//assign v_3[116] = {16'd0, decom_out[116] + v_in_3[116] + e2_ext[116]};
//assign v_3[117] = {16'd0, decom_out[117] + v_in_3[117] + e2_ext[117]};
//assign v_3[118] = {16'd0, decom_out[118] + v_in_3[118] + e2_ext[118]};
//assign v_3[119] = {16'd0, decom_out[119] + v_in_3[119] + e2_ext[119]};
//assign v_3[120] = {16'd0, decom_out[120] + v_in_3[120] + e2_ext[120]};
//assign v_3[121] = {16'd0, decom_out[121] + v_in_3[121] + e2_ext[121]};
//assign v_3[122] = {16'd0, decom_out[122] + v_in_3[122] + e2_ext[122]};
//assign v_3[123] = {16'd0, decom_out[123] + v_in_3[123] + e2_ext[123]};
//assign v_3[124] = {16'd0, decom_out[124] + v_in_3[124] + e2_ext[124]};
//assign v_3[125] = {16'd0, decom_out[125] + v_in_3[125] + e2_ext[125]};
//assign v_3[126] = {16'd0, decom_out[126] + v_in_3[126] + e2_ext[126]};
//assign v_3[127] = {16'd0, decom_out[127] + v_in_3[127] + e2_ext[127]};
//assign v_3[128] = {16'd0, decom_out[128] + v_in_3[128] + e2_ext[128]};
//assign v_3[129] = {16'd0, decom_out[129] + v_in_3[129] + e2_ext[129]};
//assign v_3[130] = {16'd0, decom_out[130] + v_in_3[130] + e2_ext[130]};
//assign v_3[131] = {16'd0, decom_out[131] + v_in_3[131] + e2_ext[131]};
//assign v_3[132] = {16'd0, decom_out[132] + v_in_3[132] + e2_ext[132]};
//assign v_3[133] = {16'd0, decom_out[133] + v_in_3[133] + e2_ext[133]};
//assign v_3[134] = {16'd0, decom_out[134] + v_in_3[134] + e2_ext[134]};
//assign v_3[135] = {16'd0, decom_out[135] + v_in_3[135] + e2_ext[135]};
//assign v_3[136] = {16'd0, decom_out[136] + v_in_3[136] + e2_ext[136]};
//assign v_3[137] = {16'd0, decom_out[137] + v_in_3[137] + e2_ext[137]};
//assign v_3[138] = {16'd0, decom_out[138] + v_in_3[138] + e2_ext[138]};
//assign v_3[139] = {16'd0, decom_out[139] + v_in_3[139] + e2_ext[139]};
//assign v_3[140] = {16'd0, decom_out[140] + v_in_3[140] + e2_ext[140]};
//assign v_3[141] = {16'd0, decom_out[141] + v_in_3[141] + e2_ext[141]};
//assign v_3[142] = {16'd0, decom_out[142] + v_in_3[142] + e2_ext[142]};
//assign v_3[143] = {16'd0, decom_out[143] + v_in_3[143] + e2_ext[143]};
//assign v_3[144] = {16'd0, decom_out[144] + v_in_3[144] + e2_ext[144]};
//assign v_3[145] = {16'd0, decom_out[145] + v_in_3[145] + e2_ext[145]};
//assign v_3[146] = {16'd0, decom_out[146] + v_in_3[146] + e2_ext[146]};
//assign v_3[147] = {16'd0, decom_out[147] + v_in_3[147] + e2_ext[147]};
//assign v_3[148] = {16'd0, decom_out[148] + v_in_3[148] + e2_ext[148]};
//assign v_3[149] = {16'd0, decom_out[149] + v_in_3[149] + e2_ext[149]};
//assign v_3[150] = {16'd0, decom_out[150] + v_in_3[150] + e2_ext[150]};
//assign v_3[151] = {16'd0, decom_out[151] + v_in_3[151] + e2_ext[151]};
//assign v_3[152] = {16'd0, decom_out[152] + v_in_3[152] + e2_ext[152]};
//assign v_3[153] = {16'd0, decom_out[153] + v_in_3[153] + e2_ext[153]};
//assign v_3[154] = {16'd0, decom_out[154] + v_in_3[154] + e2_ext[154]};
//assign v_3[155] = {16'd0, decom_out[155] + v_in_3[155] + e2_ext[155]};
//assign v_3[156] = {16'd0, decom_out[156] + v_in_3[156] + e2_ext[156]};
//assign v_3[157] = {16'd0, decom_out[157] + v_in_3[157] + e2_ext[157]};
//assign v_3[158] = {16'd0, decom_out[158] + v_in_3[158] + e2_ext[158]};
//assign v_3[159] = {16'd0, decom_out[159] + v_in_3[159] + e2_ext[159]};
//assign v_3[160] = {16'd0, decom_out[160] + v_in_3[160] + e2_ext[160]};
//assign v_3[161] = {16'd0, decom_out[161] + v_in_3[161] + e2_ext[161]};
//assign v_3[162] = {16'd0, decom_out[162] + v_in_3[162] + e2_ext[162]};
//assign v_3[163] = {16'd0, decom_out[163] + v_in_3[163] + e2_ext[163]};
//assign v_3[164] = {16'd0, decom_out[164] + v_in_3[164] + e2_ext[164]};
//assign v_3[165] = {16'd0, decom_out[165] + v_in_3[165] + e2_ext[165]};
//assign v_3[166] = {16'd0, decom_out[166] + v_in_3[166] + e2_ext[166]};
//assign v_3[167] = {16'd0, decom_out[167] + v_in_3[167] + e2_ext[167]};
//assign v_3[168] = {16'd0, decom_out[168] + v_in_3[168] + e2_ext[168]};
//assign v_3[169] = {16'd0, decom_out[169] + v_in_3[169] + e2_ext[169]};
//assign v_3[170] = {16'd0, decom_out[170] + v_in_3[170] + e2_ext[170]};
//assign v_3[171] = {16'd0, decom_out[171] + v_in_3[171] + e2_ext[171]};
//assign v_3[172] = {16'd0, decom_out[172] + v_in_3[172] + e2_ext[172]};
//assign v_3[173] = {16'd0, decom_out[173] + v_in_3[173] + e2_ext[173]};
//assign v_3[174] = {16'd0, decom_out[174] + v_in_3[174] + e2_ext[174]};
//assign v_3[175] = {16'd0, decom_out[175] + v_in_3[175] + e2_ext[175]};
//assign v_3[176] = {16'd0, decom_out[176] + v_in_3[176] + e2_ext[176]};
//assign v_3[177] = {16'd0, decom_out[177] + v_in_3[177] + e2_ext[177]};
//assign v_3[178] = {16'd0, decom_out[178] + v_in_3[178] + e2_ext[178]};
//assign v_3[179] = {16'd0, decom_out[179] + v_in_3[179] + e2_ext[179]};
//assign v_3[180] = {16'd0, decom_out[180] + v_in_3[180] + e2_ext[180]};
//assign v_3[181] = {16'd0, decom_out[181] + v_in_3[181] + e2_ext[181]};
//assign v_3[182] = {16'd0, decom_out[182] + v_in_3[182] + e2_ext[182]};
//assign v_3[183] = {16'd0, decom_out[183] + v_in_3[183] + e2_ext[183]};
//assign v_3[184] = {16'd0, decom_out[184] + v_in_3[184] + e2_ext[184]};
//assign v_3[185] = {16'd0, decom_out[185] + v_in_3[185] + e2_ext[185]};
//assign v_3[186] = {16'd0, decom_out[186] + v_in_3[186] + e2_ext[186]};
//assign v_3[187] = {16'd0, decom_out[187] + v_in_3[187] + e2_ext[187]};
//assign v_3[188] = {16'd0, decom_out[188] + v_in_3[188] + e2_ext[188]};
//assign v_3[189] = {16'd0, decom_out[189] + v_in_3[189] + e2_ext[189]};
//assign v_3[190] = {16'd0, decom_out[190] + v_in_3[190] + e2_ext[190]};
//assign v_3[191] = {16'd0, decom_out[191] + v_in_3[191] + e2_ext[191]};
//assign v_3[192] = {16'd0, decom_out[192] + v_in_3[192] + e2_ext[192]};
//assign v_3[193] = {16'd0, decom_out[193] + v_in_3[193] + e2_ext[193]};
//assign v_3[194] = {16'd0, decom_out[194] + v_in_3[194] + e2_ext[194]};
//assign v_3[195] = {16'd0, decom_out[195] + v_in_3[195] + e2_ext[195]};
//assign v_3[196] = {16'd0, decom_out[196] + v_in_3[196] + e2_ext[196]};
//assign v_3[197] = {16'd0, decom_out[197] + v_in_3[197] + e2_ext[197]};
//assign v_3[198] = {16'd0, decom_out[198] + v_in_3[198] + e2_ext[198]};
//assign v_3[199] = {16'd0, decom_out[199] + v_in_3[199] + e2_ext[199]};
//assign v_3[200] = {16'd0, decom_out[200] + v_in_3[200] + e2_ext[200]};
//assign v_3[201] = {16'd0, decom_out[201] + v_in_3[201] + e2_ext[201]};
//assign v_3[202] = {16'd0, decom_out[202] + v_in_3[202] + e2_ext[202]};
//assign v_3[203] = {16'd0, decom_out[203] + v_in_3[203] + e2_ext[203]};
//assign v_3[204] = {16'd0, decom_out[204] + v_in_3[204] + e2_ext[204]};
//assign v_3[205] = {16'd0, decom_out[205] + v_in_3[205] + e2_ext[205]};
//assign v_3[206] = {16'd0, decom_out[206] + v_in_3[206] + e2_ext[206]};
//assign v_3[207] = {16'd0, decom_out[207] + v_in_3[207] + e2_ext[207]};
//assign v_3[208] = {16'd0, decom_out[208] + v_in_3[208] + e2_ext[208]};
//assign v_3[209] = {16'd0, decom_out[209] + v_in_3[209] + e2_ext[209]};
//assign v_3[210] = {16'd0, decom_out[210] + v_in_3[210] + e2_ext[210]};
//assign v_3[211] = {16'd0, decom_out[211] + v_in_3[211] + e2_ext[211]};
//assign v_3[212] = {16'd0, decom_out[212] + v_in_3[212] + e2_ext[212]};
//assign v_3[213] = {16'd0, decom_out[213] + v_in_3[213] + e2_ext[213]};
//assign v_3[214] = {16'd0, decom_out[214] + v_in_3[214] + e2_ext[214]};
//assign v_3[215] = {16'd0, decom_out[215] + v_in_3[215] + e2_ext[215]};
//assign v_3[216] = {16'd0, decom_out[216] + v_in_3[216] + e2_ext[216]};
//assign v_3[217] = {16'd0, decom_out[217] + v_in_3[217] + e2_ext[217]};
//assign v_3[218] = {16'd0, decom_out[218] + v_in_3[218] + e2_ext[218]};
//assign v_3[219] = {16'd0, decom_out[219] + v_in_3[219] + e2_ext[219]};
//assign v_3[220] = {16'd0, decom_out[220] + v_in_3[220] + e2_ext[220]};
//assign v_3[221] = {16'd0, decom_out[221] + v_in_3[221] + e2_ext[221]};
//assign v_3[222] = {16'd0, decom_out[222] + v_in_3[222] + e2_ext[222]};
//assign v_3[223] = {16'd0, decom_out[223] + v_in_3[223] + e2_ext[223]};
//assign v_3[224] = {16'd0, decom_out[224] + v_in_3[224] + e2_ext[224]};
//assign v_3[225] = {16'd0, decom_out[225] + v_in_3[225] + e2_ext[225]};
//assign v_3[226] = {16'd0, decom_out[226] + v_in_3[226] + e2_ext[226]};
//assign v_3[227] = {16'd0, decom_out[227] + v_in_3[227] + e2_ext[227]};
//assign v_3[228] = {16'd0, decom_out[228] + v_in_3[228] + e2_ext[228]};
//assign v_3[229] = {16'd0, decom_out[229] + v_in_3[229] + e2_ext[229]};
//assign v_3[230] = {16'd0, decom_out[230] + v_in_3[230] + e2_ext[230]};
//assign v_3[231] = {16'd0, decom_out[231] + v_in_3[231] + e2_ext[231]};
//assign v_3[232] = {16'd0, decom_out[232] + v_in_3[232] + e2_ext[232]};
//assign v_3[233] = {16'd0, decom_out[233] + v_in_3[233] + e2_ext[233]};
//assign v_3[234] = {16'd0, decom_out[234] + v_in_3[234] + e2_ext[234]};
//assign v_3[235] = {16'd0, decom_out[235] + v_in_3[235] + e2_ext[235]};
//assign v_3[236] = {16'd0, decom_out[236] + v_in_3[236] + e2_ext[236]};
//assign v_3[237] = {16'd0, decom_out[237] + v_in_3[237] + e2_ext[237]};
//assign v_3[238] = {16'd0, decom_out[238] + v_in_3[238] + e2_ext[238]};
//assign v_3[239] = {16'd0, decom_out[239] + v_in_3[239] + e2_ext[239]};
//assign v_3[240] = {16'd0, decom_out[240] + v_in_3[240] + e2_ext[240]};
//assign v_3[241] = {16'd0, decom_out[241] + v_in_3[241] + e2_ext[241]};
//assign v_3[242] = {16'd0, decom_out[242] + v_in_3[242] + e2_ext[242]};
//assign v_3[243] = {16'd0, decom_out[243] + v_in_3[243] + e2_ext[243]};
//assign v_3[244] = {16'd0, decom_out[244] + v_in_3[244] + e2_ext[244]};
//assign v_3[245] = {16'd0, decom_out[245] + v_in_3[245] + e2_ext[245]};
//assign v_3[246] = {16'd0, decom_out[246] + v_in_3[246] + e2_ext[246]};
//assign v_3[247] = {16'd0, decom_out[247] + v_in_3[247] + e2_ext[247]};
//assign v_3[248] = {16'd0, decom_out[248] + v_in_3[248] + e2_ext[248]};
//assign v_3[249] = {16'd0, decom_out[249] + v_in_3[249] + e2_ext[249]};
//assign v_3[250] = {16'd0, decom_out[250] + v_in_3[250] + e2_ext[250]};
//assign v_3[251] = {16'd0, decom_out[251] + v_in_3[251] + e2_ext[251]};
//assign v_3[252] = {16'd0, decom_out[252] + v_in_3[252] + e2_ext[252]};
//assign v_3[253] = {16'd0, decom_out[253] + v_in_3[253] + e2_ext[253]};
//assign v_3[254] = {16'd0, decom_out[254] + v_in_3[254] + e2_ext[254]};
//assign v_3[255] = {16'd0, decom_out[255] + v_in_3[255] + e2_ext[255]};

 
//compress_module compress_1 (
//    .x(16),
//    .d(u_1[0]),
//    .result(com_out[0])
//);

//compress_module compress_2 (
//    .x(16),
//    .d(u_1[1]),
//    .result(com_out[1])
//);

//compress_module compress_3 (
//    .x(16),
//    .d(u_1[2]),
//    .result(com_out[2])
//);

//compress_module compress_4 (
//    .x(16),
//    .d(u_1[3]),
//    .result(com_out[3])
//);

//compress_module compress_5 (
//    .x(16),
//    .d(u_1[4]),
//    .result(com_out[4])
//);

//compress_module compress_6 (
//    .x(16),
//    .d(u_1[5]),
//    .result(com_out[5])
//);

//compress_module compress_7 (
//    .x(16),
//    .d(u_1[6]),
//    .result(com_out[6])
//);

//compress_module compress_8 (
//    .x(16),
//    .d(u_1[7]),
//    .result(com_out[7])
//);

//compress_module compress_9 (
//    .x(16),
//    .d(u_1[8]),
//    .result(com_out[8])
//);

//compress_module compress_10 (
//    .x(16),
//    .d(u_1[9]),
//    .result(com_out[9])
//);

//compress_module compress_11 (
//    .x(16),
//    .d(u_1[10]),
//    .result(com_out[10])
//);

//compress_module compress_12 (
//    .x(16),
//    .d(u_1[11]),
//    .result(com_out[11])
//);

//compress_module compress_13 (
//    .x(16),
//    .d(u_1[12]),
//    .result(com_out[12])
//);

//compress_module compress_14 (
//    .x(16),
//    .d(u_1[13]),
//    .result(com_out[13])
//);

//compress_module compress_15 (
//    .x(16),
//    .d(u_1[14]),
//    .result(com_out[14])
//);

//compress_module compress_16 (
//    .x(16),
//    .d(u_1[15]),
//    .result(com_out[15])
//);

//compress_module compress_17 (
//    .x(16),
//    .d(u_1[16]),
//    .result(com_out[16])
//);

//compress_module compress_18 (
//    .x(16),
//    .d(u_1[17]),
//    .result(com_out[17])
//);

//compress_module compress_19 (
//    .x(16),
//    .d(u_1[18]),
//    .result(com_out[18])
//);

//compress_module compress_20 (
//    .x(16),
//    .d(u_1[19]),
//    .result(com_out[19])
//);

//compress_module compress_21 (
//    .x(16),
//    .d(u_1[20]),
//    .result(com_out[20])
//);

//compress_module compress_22 (
//    .x(16),
//    .d(u_1[21]),
//    .result(com_out[21])
//);

//compress_module compress_23 (
//    .x(16),
//    .d(u_1[22]),
//    .result(com_out[22])
//);

//compress_module compress_24 (
//    .x(16),
//    .d(u_1[23]),
//    .result(com_out[23])
//);

//compress_module compress_25 (
//    .x(16),
//    .d(u_1[24]),
//    .result(com_out[24])
//);

//compress_module compress_26 (
//    .x(16),
//    .d(u_1[25]),
//    .result(com_out[25])
//);

//compress_module compress_27 (
//    .x(16),
//    .d(u_1[26]),
//    .result(com_out[26])
//);

//compress_module compress_28 (
//    .x(16),
//    .d(u_1[27]),
//    .result(com_out[27])
//);

//compress_module compress_29 (
//    .x(16),
//    .d(u_1[28]),
//    .result(com_out[28])
//);

//compress_module compress_30 (
//    .x(16),
//    .d(u_1[29]),
//    .result(com_out[29])
//);

//compress_module compress_31 (
//    .x(16),
//    .d(u_1[30]),
//    .result(com_out[30])
//);

//compress_module compress_32 (
//    .x(16),
//    .d(u_1[31]),
//    .result(com_out[31])
//);

//compress_module compress_33 (
//    .x(16),
//    .d(u_1[32]),
//    .result(com_out[32])
//);

//compress_module compress_34 (
//    .x(16),
//    .d(u_1[33]),
//    .result(com_out[33])
//);

//compress_module compress_35 (
//    .x(16),
//    .d(u_1[34]),
//    .result(com_out[34])
//);

//compress_module compress_36 (
//    .x(16),
//    .d(u_1[35]),
//    .result(com_out[35])
//);

//compress_module compress_37 (
//    .x(16),
//    .d(u_1[36]),
//    .result(com_out[36])
//);

//compress_module compress_38 (
//    .x(16),
//    .d(u_1[37]),
//    .result(com_out[37])
//);

//compress_module compress_39 (
//    .x(16),
//    .d(u_1[38]),
//    .result(com_out[38])
//);

//compress_module compress_40 (
//    .x(16),
//    .d(u_1[39]),
//    .result(com_out[39])
//);

//compress_module compress_41 (
//    .x(16),
//    .d(u_1[40]),
//    .result(com_out[40])
//);

//compress_module compress_42 (
//    .x(16),
//    .d(u_1[41]),
//    .result(com_out[41])
//);

//compress_module compress_43 (
//    .x(16),
//    .d(u_1[42]),
//    .result(com_out[42])
//);

//compress_module compress_44 (
//    .x(16),
//    .d(u_1[43]),
//    .result(com_out[43])
//);

//compress_module compress_45 (
//    .x(16),
//    .d(u_1[44]),
//    .result(com_out[44])
//);

//compress_module compress_46 (
//    .x(16),
//    .d(u_1[45]),
//    .result(com_out[45])
//);

//compress_module compress_47 (
//    .x(16),
//    .d(u_1[46]),
//    .result(com_out[46])
//);

//compress_module compress_48 (
//    .x(16),
//    .d(u_1[47]),
//    .result(com_out[47])
//);

//compress_module compress_49 (
//    .x(16),
//    .d(u_1[48]),
//    .result(com_out[48])
//);

//compress_module compress_50 (
//    .x(16),
//    .d(u_1[49]),
//    .result(com_out[49])
//);

//compress_module compress_51 (
//    .x(16),
//    .d(u_1[50]),
//    .result(com_out[50])
//);

//compress_module compress_52 (
//    .x(16),
//    .d(u_1[51]),
//    .result(com_out[51])
//);

//compress_module compress_53 (
//    .x(16),
//    .d(u_1[52]),
//    .result(com_out[52])
//);

//compress_module compress_54 (
//    .x(16),
//    .d(u_1[53]),
//    .result(com_out[53])
//);

//compress_module compress_55 (
//    .x(16),
//    .d(u_1[54]),
//    .result(com_out[54])
//);

//compress_module compress_56 (
//    .x(16),
//    .d(u_1[55]),
//    .result(com_out[55])
//);

//compress_module compress_57 (
//    .x(16),
//    .d(u_1[56]),
//    .result(com_out[56])
//);

//compress_module compress_58 (
//    .x(16),
//    .d(u_1[57]),
//    .result(com_out[57])
//);

//compress_module compress_59 (
//    .x(16),
//    .d(u_1[58]),
//    .result(com_out[58])
//);

//compress_module compress_60 (
//    .x(16),
//    .d(u_1[59]),
//    .result(com_out[59])
//);

//compress_module compress_61 (
//    .x(16),
//    .d(u_1[60]),
//    .result(com_out[60])
//);

//compress_module compress_62 (
//    .x(16),
//    .d(u_1[61]),
//    .result(com_out[61])
//);

//compress_module compress_63 (
//    .x(16),
//    .d(u_1[62]),
//    .result(com_out[62])
//);

//compress_module compress_64 (
//    .x(16),
//    .d(u_1[63]),
//    .result(com_out[63])
//);

//compress_module compress_65 (
//    .x(16),
//    .d(u_1[64]),
//    .result(com_out[64])
//);

//compress_module compress_66 (
//    .x(16),
//    .d(u_1[65]),
//    .result(com_out[65])
//);

//compress_module compress_67 (
//    .x(16),
//    .d(u_1[66]),
//    .result(com_out[66])
//);

//compress_module compress_68 (
//    .x(16),
//    .d(u_1[67]),
//    .result(com_out[67])
//);

//compress_module compress_69 (
//    .x(16),
//    .d(u_1[68]),
//    .result(com_out[68])
//);

//compress_module compress_70 (
//    .x(16),
//    .d(u_1[69]),
//    .result(com_out[69])
//);

//compress_module compress_71 (
//    .x(16),
//    .d(u_1[70]),
//    .result(com_out[70])
//);

//compress_module compress_72 (
//    .x(16),
//    .d(u_1[71]),
//    .result(com_out[71])
//);

//compress_module compress_73 (
//    .x(16),
//    .d(u_1[72]),
//    .result(com_out[72])
//);

//compress_module compress_74 (
//    .x(16),
//    .d(u_1[73]),
//    .result(com_out[73])
//);

//compress_module compress_75 (
//    .x(16),
//    .d(u_1[74]),
//    .result(com_out[74])
//);

//compress_module compress_76 (
//    .x(16),
//    .d(u_1[75]),
//    .result(com_out[75])
//);

//compress_module compress_77 (
//    .x(16),
//    .d(u_1[76]),
//    .result(com_out[76])
//);

//compress_module compress_78 (
//    .x(16),
//    .d(u_1[77]),
//    .result(com_out[77])
//);

//compress_module compress_79 (
//    .x(16),
//    .d(u_1[78]),
//    .result(com_out[78])
//);

//compress_module compress_80 (
//    .x(16),
//    .d(u_1[79]),
//    .result(com_out[79])
//);

//compress_module compress_81 (
//    .x(16),
//    .d(u_1[80]),
//    .result(com_out[80])
//);

//compress_module compress_82 (
//    .x(16),
//    .d(u_1[81]),
//    .result(com_out[81])
//);

//compress_module compress_83 (
//    .x(16),
//    .d(u_1[82]),
//    .result(com_out[82])
//);

//compress_module compress_84 (
//    .x(16),
//    .d(u_1[83]),
//    .result(com_out[83])
//);

//compress_module compress_85 (
//    .x(16),
//    .d(u_1[84]),
//    .result(com_out[84])
//);

//compress_module compress_86 (
//    .x(16),
//    .d(u_1[85]),
//    .result(com_out[85])
//);

//compress_module compress_87 (
//    .x(16),
//    .d(u_1[86]),
//    .result(com_out[86])
//);

//compress_module compress_88 (
//    .x(16),
//    .d(u_1[87]),
//    .result(com_out[87])
//);

//compress_module compress_89 (
//    .x(16),
//    .d(u_1[88]),
//    .result(com_out[88])
//);

//compress_module compress_90 (
//    .x(16),
//    .d(u_1[89]),
//    .result(com_out[89])
//);

//compress_module compress_91 (
//    .x(16),
//    .d(u_1[90]),
//    .result(com_out[90])
//);

//compress_module compress_92 (
//    .x(16),
//    .d(u_1[91]),
//    .result(com_out[91])
//);

//compress_module compress_93 (
//    .x(16),
//    .d(u_1[92]),
//    .result(com_out[92])
//);

//compress_module compress_94 (
//    .x(16),
//    .d(u_1[93]),
//    .result(com_out[93])
//);

//compress_module compress_95 (
//    .x(16),
//    .d(u_1[94]),
//    .result(com_out[94])
//);

//compress_module compress_96 (
//    .x(16),
//    .d(u_1[95]),
//    .result(com_out[95])
//);

//compress_module compress_97 (
//    .x(16),
//    .d(u_1[96]),
//    .result(com_out[96])
//);

//compress_module compress_98 (
//    .x(16),
//    .d(u_1[97]),
//    .result(com_out[97])
//);

//compress_module compress_99 (
//    .x(16),
//    .d(u_1[98]),
//    .result(com_out[98])
//);

//compress_module compress_100 (
//    .x(16),
//    .d(u_1[99]),
//    .result(com_out[99])
//);

//compress_module compress_101 (
//    .x(16),
//    .d(u_1[100]),
//    .result(com_out[100])
//);

//compress_module compress_102 (
//    .x(16),
//    .d(u_1[101]),
//    .result(com_out[101])
//);

//compress_module compress_103 (
//    .x(16),
//    .d(u_1[102]),
//    .result(com_out[102])
//);

//compress_module compress_104 (
//    .x(16),
//    .d(u_1[103]),
//    .result(com_out[103])
//);

//compress_module compress_105 (
//    .x(16),
//    .d(u_1[104]),
//    .result(com_out[104])
//);

//compress_module compress_106 (
//    .x(16),
//    .d(u_1[105]),
//    .result(com_out[105])
//);

//compress_module compress_107 (
//    .x(16),
//    .d(u_1[106]),
//    .result(com_out[106])
//);

//compress_module compress_108 (
//    .x(16),
//    .d(u_1[107]),
//    .result(com_out[107])
//);

//compress_module compress_109 (
//    .x(16),
//    .d(u_1[108]),
//    .result(com_out[108])
//);

//compress_module compress_110 (
//    .x(16),
//    .d(u_1[109]),
//    .result(com_out[109])
//);

//compress_module compress_111 (
//    .x(16),
//    .d(u_1[110]),
//    .result(com_out[110])
//);

//compress_module compress_112 (
//    .x(16),
//    .d(u_1[111]),
//    .result(com_out[111])
//);

//compress_module compress_113 (
//    .x(16),
//    .d(u_1[112]),
//    .result(com_out[112])
//);

//compress_module compress_114 (
//    .x(16),
//    .d(u_1[113]),
//    .result(com_out[113])
//);

//compress_module compress_115 (
//    .x(16),
//    .d(u_1[114]),
//    .result(com_out[114])
//);

//compress_module compress_116 (
//    .x(16),
//    .d(u_1[115]),
//    .result(com_out[115])
//);

//compress_module compress_117 (
//    .x(16),
//    .d(u_1[116]),
//    .result(com_out[116])
//);

//compress_module compress_118 (
//    .x(16),
//    .d(u_1[117]),
//    .result(com_out[117])
//);

//compress_module compress_119 (
//    .x(16),
//    .d(u_1[118]),
//    .result(com_out[118])
//);

//compress_module compress_120 (
//    .x(16),
//    .d(u_1[119]),
//    .result(com_out[119])
//);

//compress_module compress_121 (
//    .x(16),
//    .d(u_1[120]),
//    .result(com_out[120])
//);

//compress_module compress_122 (
//    .x(16),
//    .d(u_1[121]),
//    .result(com_out[121])
//);

//compress_module compress_123 (
//    .x(16),
//    .d(u_1[122]),
//    .result(com_out[122])
//);

//compress_module compress_124 (
//    .x(16),
//    .d(u_1[123]),
//    .result(com_out[123])
//);

//compress_module compress_125 (
//    .x(16),
//    .d(u_1[124]),
//    .result(com_out[124])
//);

//compress_module compress_126 (
//    .x(16),
//    .d(u_1[125]),
//    .result(com_out[125])
//);

//compress_module compress_127 (
//    .x(16),
//    .d(u_1[126]),
//    .result(com_out[126])
//);

//compress_module compress_128 (
//    .x(16),
//    .d(u_1[127]),
//    .result(com_out[127])
//);

//compress_module compress_129 (
//    .x(16),
//    .d(u_1[128]),
//    .result(com_out[128])
//);

//compress_module compress_130 (
//    .x(16),
//    .d(u_1[129]),
//    .result(com_out[129])
//);

//compress_module compress_131 (
//    .x(16),
//    .d(u_1[130]),
//    .result(com_out[130])
//);

//compress_module compress_132 (
//    .x(16),
//    .d(u_1[131]),
//    .result(com_out[131])
//);

//compress_module compress_133 (
//    .x(16),
//    .d(u_1[132]),
//    .result(com_out[132])
//);

//compress_module compress_134 (
//    .x(16),
//    .d(u_1[133]),
//    .result(com_out[133])
//);

//compress_module compress_135 (
//    .x(16),
//    .d(u_1[134]),
//    .result(com_out[134])
//);

//compress_module compress_136 (
//    .x(16),
//    .d(u_1[135]),
//    .result(com_out[135])
//);

//compress_module compress_137 (
//    .x(16),
//    .d(u_1[136]),
//    .result(com_out[136])
//);

//compress_module compress_138 (
//    .x(16),
//    .d(u_1[137]),
//    .result(com_out[137])
//);

//compress_module compress_139 (
//    .x(16),
//    .d(u_1[138]),
//    .result(com_out[138])
//);

//compress_module compress_140 (
//    .x(16),
//    .d(u_1[139]),
//    .result(com_out[139])
//);

//compress_module compress_141 (
//    .x(16),
//    .d(u_1[140]),
//    .result(com_out[140])
//);

//compress_module compress_142 (
//    .x(16),
//    .d(u_1[141]),
//    .result(com_out[141])
//);

//compress_module compress_143 (
//    .x(16),
//    .d(u_1[142]),
//    .result(com_out[142])
//);

//compress_module compress_144 (
//    .x(16),
//    .d(u_1[143]),
//    .result(com_out[143])
//);

//compress_module compress_145 (
//    .x(16),
//    .d(u_1[144]),
//    .result(com_out[144])
//);

//compress_module compress_146 (
//    .x(16),
//    .d(u_1[145]),
//    .result(com_out[145])
//);

//compress_module compress_147 (
//    .x(16),
//    .d(u_1[146]),
//    .result(com_out[146])
//);

//compress_module compress_148 (
//    .x(16),
//    .d(u_1[147]),
//    .result(com_out[147])
//);

//compress_module compress_149 (
//    .x(16),
//    .d(u_1[148]),
//    .result(com_out[148])
//);

//compress_module compress_150 (
//    .x(16),
//    .d(u_1[149]),
//    .result(com_out[149])
//);

//compress_module compress_151 (
//    .x(16),
//    .d(u_1[150]),
//    .result(com_out[150])
//);

//compress_module compress_152 (
//    .x(16),
//    .d(u_1[151]),
//    .result(com_out[151])
//);

//compress_module compress_153 (
//    .x(16),
//    .d(u_1[152]),
//    .result(com_out[152])
//);

//compress_module compress_154 (
//    .x(16),
//    .d(u_1[153]),
//    .result(com_out[153])
//);

//compress_module compress_155 (
//    .x(16),
//    .d(u_1[154]),
//    .result(com_out[154])
//);

//compress_module compress_156 (
//    .x(16),
//    .d(u_1[155]),
//    .result(com_out[155])
//);

//compress_module compress_157 (
//    .x(16),
//    .d(u_1[156]),
//    .result(com_out[156])
//);

//compress_module compress_158 (
//    .x(16),
//    .d(u_1[157]),
//    .result(com_out[157])
//);

//compress_module compress_159 (
//    .x(16),
//    .d(u_1[158]),
//    .result(com_out[158])
//);

//compress_module compress_160 (
//    .x(16),
//    .d(u_1[159]),
//    .result(com_out[159])
//);

//compress_module compress_161 (
//    .x(16),
//    .d(u_1[160]),
//    .result(com_out[160])
//);

//compress_module compress_162 (
//    .x(16),
//    .d(u_1[161]),
//    .result(com_out[161])
//);

//compress_module compress_163 (
//    .x(16),
//    .d(u_1[162]),
//    .result(com_out[162])
//);

//compress_module compress_164 (
//    .x(16),
//    .d(u_1[163]),
//    .result(com_out[163])
//);

//compress_module compress_165 (
//    .x(16),
//    .d(u_1[164]),
//    .result(com_out[164])
//);

//compress_module compress_166 (
//    .x(16),
//    .d(u_1[165]),
//    .result(com_out[165])
//);

//compress_module compress_167 (
//    .x(16),
//    .d(u_1[166]),
//    .result(com_out[166])
//);

//compress_module compress_168 (
//    .x(16),
//    .d(u_1[167]),
//    .result(com_out[167])
//);

//compress_module compress_169 (
//    .x(16),
//    .d(u_1[168]),
//    .result(com_out[168])
//);

//compress_module compress_170 (
//    .x(16),
//    .d(u_1[169]),
//    .result(com_out[169])
//);

//compress_module compress_171 (
//    .x(16),
//    .d(u_1[170]),
//    .result(com_out[170])
//);

//compress_module compress_172 (
//    .x(16),
//    .d(u_1[171]),
//    .result(com_out[171])
//);

//compress_module compress_173 (
//    .x(16),
//    .d(u_1[172]),
//    .result(com_out[172])
//);

//compress_module compress_174 (
//    .x(16),
//    .d(u_1[173]),
//    .result(com_out[173])
//);

//compress_module compress_175 (
//    .x(16),
//    .d(u_1[174]),
//    .result(com_out[174])
//);

//compress_module compress_176 (
//    .x(16),
//    .d(u_1[175]),
//    .result(com_out[175])
//);

//compress_module compress_177 (
//    .x(16),
//    .d(u_1[176]),
//    .result(com_out[176])
//);

//compress_module compress_178 (
//    .x(16),
//    .d(u_1[177]),
//    .result(com_out[177])
//);

//compress_module compress_179 (
//    .x(16),
//    .d(u_1[178]),
//    .result(com_out[178])
//);

//compress_module compress_180 (
//    .x(16),
//    .d(u_1[179]),
//    .result(com_out[179])
//);

//compress_module compress_181 (
//    .x(16),
//    .d(u_1[180]),
//    .result(com_out[180])
//);

//compress_module compress_182 (
//    .x(16),
//    .d(u_1[181]),
//    .result(com_out[181])
//);

//compress_module compress_183 (
//    .x(16),
//    .d(u_1[182]),
//    .result(com_out[182])
//);

//compress_module compress_184 (
//    .x(16),
//    .d(u_1[183]),
//    .result(com_out[183])
//);

//compress_module compress_185 (
//    .x(16),
//    .d(u_1[184]),
//    .result(com_out[184])
//);

//compress_module compress_186 (
//    .x(16),
//    .d(u_1[185]),
//    .result(com_out[185])
//);

//compress_module compress_187 (
//    .x(16),
//    .d(u_1[186]),
//    .result(com_out[186])
//);

//compress_module compress_188 (
//    .x(16),
//    .d(u_1[187]),
//    .result(com_out[187])
//);

//compress_module compress_189 (
//    .x(16),
//    .d(u_1[188]),
//    .result(com_out[188])
//);

//compress_module compress_190 (
//    .x(16),
//    .d(u_1[189]),
//    .result(com_out[189])
//);

//compress_module compress_191 (
//    .x(16),
//    .d(u_1[190]),
//    .result(com_out[190])
//);

//compress_module compress_192 (
//    .x(16),
//    .d(u_1[191]),
//    .result(com_out[191])
//);

//compress_module compress_193 (
//    .x(16),
//    .d(u_1[192]),
//    .result(com_out[192])
//);

//compress_module compress_194 (
//    .x(16),
//    .d(u_1[193]),
//    .result(com_out[193])
//);

//compress_module compress_195 (
//    .x(16),
//    .d(u_1[194]),
//    .result(com_out[194])
//);

//compress_module compress_196 (
//    .x(16),
//    .d(u_1[195]),
//    .result(com_out[195])
//);

//compress_module compress_197 (
//    .x(16),
//    .d(u_1[196]),
//    .result(com_out[196])
//);

//compress_module compress_198 (
//    .x(16),
//    .d(u_1[197]),
//    .result(com_out[197])
//);

//compress_module compress_199 (
//    .x(16),
//    .d(u_1[198]),
//    .result(com_out[198])
//);

//compress_module compress_200 (
//    .x(16),
//    .d(u_1[199]),
//    .result(com_out[199])
//);

//compress_module compress_201 (
//    .x(16),
//    .d(u_1[200]),
//    .result(com_out[200])
//);

//compress_module compress_202 (
//    .x(16),
//    .d(u_1[201]),
//    .result(com_out[201])
//);

//compress_module compress_203 (
//    .x(16),
//    .d(u_1[202]),
//    .result(com_out[202])
//);

//compress_module compress_204 (
//    .x(16),
//    .d(u_1[203]),
//    .result(com_out[203])
//);

//compress_module compress_205 (
//    .x(16),
//    .d(u_1[204]),
//    .result(com_out[204])
//);

//compress_module compress_206 (
//    .x(16),
//    .d(u_1[205]),
//    .result(com_out[205])
//);

//compress_module compress_207 (
//    .x(16),
//    .d(u_1[206]),
//    .result(com_out[206])
//);

//compress_module compress_208 (
//    .x(16),
//    .d(u_1[207]),
//    .result(com_out[207])
//);

//compress_module compress_209 (
//    .x(16),
//    .d(u_1[208]),
//    .result(com_out[208])
//);

//compress_module compress_210 (
//    .x(16),
//    .d(u_1[209]),
//    .result(com_out[209])
//);

//compress_module compress_211 (
//    .x(16),
//    .d(u_1[210]),
//    .result(com_out[210])
//);

//compress_module compress_212 (
//    .x(16),
//    .d(u_1[211]),
//    .result(com_out[211])
//);

//compress_module compress_213 (
//    .x(16),
//    .d(u_1[212]),
//    .result(com_out[212])
//);

//compress_module compress_214 (
//    .x(16),
//    .d(u_1[213]),
//    .result(com_out[213])
//);

//compress_module compress_215 (
//    .x(16),
//    .d(u_1[214]),
//    .result(com_out[214])
//);

//compress_module compress_216 (
//    .x(16),
//    .d(u_1[215]),
//    .result(com_out[215])
//);

//compress_module compress_217 (
//    .x(16),
//    .d(u_1[216]),
//    .result(com_out[216])
//);

//compress_module compress_218 (
//    .x(16),
//    .d(u_1[217]),
//    .result(com_out[217])
//);

//compress_module compress_219 (
//    .x(16),
//    .d(u_1[218]),
//    .result(com_out[218])
//);

//compress_module compress_220 (
//    .x(16),
//    .d(u_1[219]),
//    .result(com_out[219])
//);

//compress_module compress_221 (
//    .x(16),
//    .d(u_1[220]),
//    .result(com_out[220])
//);

//compress_module compress_222 (
//    .x(16),
//    .d(u_1[221]),
//    .result(com_out[221])
//);

//compress_module compress_223 (
//    .x(16),
//    .d(u_1[222]),
//    .result(com_out[222])
//);

//compress_module compress_224 (
//    .x(16),
//    .d(u_1[223]),
//    .result(com_out[223])
//);

//compress_module compress_225 (
//    .x(16),
//    .d(u_1[224]),
//    .result(com_out[224])
//);

//compress_module compress_226 (
//    .x(16),
//    .d(u_1[225]),
//    .result(com_out[225])
//);

//compress_module compress_227 (
//    .x(16),
//    .d(u_1[226]),
//    .result(com_out[226])
//);

//compress_module compress_228 (
//    .x(16),
//    .d(u_1[227]),
//    .result(com_out[227])
//);

//compress_module compress_229 (
//    .x(16),
//    .d(u_1[228]),
//    .result(com_out[228])
//);

//compress_module compress_230 (
//    .x(16),
//    .d(u_1[229]),
//    .result(com_out[229])
//);

//compress_module compress_231 (
//    .x(16),
//    .d(u_1[230]),
//    .result(com_out[230])
//);

//compress_module compress_232 (
//    .x(16),
//    .d(u_1[231]),
//    .result(com_out[231])
//);

//compress_module compress_233 (
//    .x(16),
//    .d(u_1[232]),
//    .result(com_out[232])
//);

//compress_module compress_234 (
//    .x(16),
//    .d(u_1[233]),
//    .result(com_out[233])
//);

//compress_module compress_235 (
//    .x(16),
//    .d(u_1[234]),
//    .result(com_out[234])
//);

//compress_module compress_236 (
//    .x(16),
//    .d(u_1[235]),
//    .result(com_out[235])
//);

//compress_module compress_237 (
//    .x(16),
//    .d(u_1[236]),
//    .result(com_out[236])
//);

//compress_module compress_238 (
//    .x(16),
//    .d(u_1[237]),
//    .result(com_out[237])
//);

//compress_module compress_239 (
//    .x(16),
//    .d(u_1[238]),
//    .result(com_out[238])
//);

//compress_module compress_240 (
//    .x(16),
//    .d(u_1[239]),
//    .result(com_out[239])
//);

//compress_module compress_241 (
//    .x(16),
//    .d(u_1[240]),
//    .result(com_out[240])
//);

//compress_module compress_242 (
//    .x(16),
//    .d(u_1[241]),
//    .result(com_out[241])
//);

//compress_module compress_243 (
//    .x(16),
//    .d(u_1[242]),
//    .result(com_out[242])
//);

//compress_module compress_244 (
//    .x(16),
//    .d(u_1[243]),
//    .result(com_out[243])
//);

//compress_module compress_245 (
//    .x(16),
//    .d(u_1[244]),
//    .result(com_out[244])
//);

//compress_module compress_246 (
//    .x(16),
//    .d(u_1[245]),
//    .result(com_out[245])
//);

//compress_module compress_247 (
//    .x(16),
//    .d(u_1[246]),
//    .result(com_out[246])
//);

//compress_module compress_248 (
//    .x(16),
//    .d(u_1[247]),
//    .result(com_out[247])
//);

//compress_module compress_249 (
//    .x(16),
//    .d(u_1[248]),
//    .result(com_out[248])
//);

//compress_module compress_250 (
//    .x(16),
//    .d(u_1[249]),
//    .result(com_out[249])
//);

//compress_module compress_251 (
//    .x(16),
//    .d(u_1[250]),
//    .result(com_out[250])
//);

//compress_module compress_252 (
//    .x(16),
//    .d(u_1[251]),
//    .result(com_out[251])
//);

//compress_module compress_253 (
//    .x(16),
//    .d(u_1[252]),
//    .result(com_out[252])
//);

//compress_module compress_254 (
//    .x(16),
//    .d(u_1[253]),
//    .result(com_out[253])
//);

//compress_module compress_255 (
//    .x(16),
//    .d(u_1[254]),
//    .result(com_out[254])
//);

//compress_module compress_256 (
//    .x(16),
//    .d(u_1[255]),
//    .result(com_out[255])
//);

//compress_module compress_257 (
//    .x(16),
//    .d(u_2[256]),
//    .result(com_out[256])
//);

//compress_module compress_258 (
//    .x(16),
//    .d(u_2[257]),
//    .result(com_out[257])
//);

//compress_module compress_259 (
//    .x(16),
//    .d(u_2[258]),
//    .result(com_out[258])
//);

//compress_module compress_260 (
//    .x(16),
//    .d(u_2[259]),
//    .result(com_out[259])
//);

//compress_module compress_261 (
//    .x(16),
//    .d(u_2[260]),
//    .result(com_out[260])
//);

//compress_module compress_262 (
//    .x(16),
//    .d(u_2[261]),
//    .result(com_out[261])
//);

//compress_module compress_263 (
//    .x(16),
//    .d(u_2[262]),
//    .result(com_out[262])
//);

//compress_module compress_264 (
//    .x(16),
//    .d(u_2[263]),
//    .result(com_out[263])
//);

//compress_module compress_265 (
//    .x(16),
//    .d(u_2[264]),
//    .result(com_out[264])
//);

//compress_module compress_266 (
//    .x(16),
//    .d(u_2[265]),
//    .result(com_out[265])
//);

//compress_module compress_267 (
//    .x(16),
//    .d(u_2[266]),
//    .result(com_out[266])
//);

//compress_module compress_268 (
//    .x(16),
//    .d(u_2[267]),
//    .result(com_out[267])
//);

//compress_module compress_269 (
//    .x(16),
//    .d(u_2[268]),
//    .result(com_out[268])
//);

//compress_module compress_270 (
//    .x(16),
//    .d(u_2[269]),
//    .result(com_out[269])
//);

//compress_module compress_271 (
//    .x(16),
//    .d(u_2[270]),
//    .result(com_out[270])
//);

//compress_module compress_272 (
//    .x(16),
//    .d(u_2[271]),
//    .result(com_out[271])
//);

//compress_module compress_273 (
//    .x(16),
//    .d(u_2[272]),
//    .result(com_out[272])
//);

//compress_module compress_274 (
//    .x(16),
//    .d(u_2[273]),
//    .result(com_out[273])
//);

//compress_module compress_275 (
//    .x(16),
//    .d(u_2[274]),
//    .result(com_out[274])
//);

//compress_module compress_276 (
//    .x(16),
//    .d(u_2[275]),
//    .result(com_out[275])
//);

//compress_module compress_277 (
//    .x(16),
//    .d(u_2[276]),
//    .result(com_out[276])
//);

//compress_module compress_278 (
//    .x(16),
//    .d(u_2[277]),
//    .result(com_out[277])
//);

//compress_module compress_279 (
//    .x(16),
//    .d(u_2[278]),
//    .result(com_out[278])
//);

//compress_module compress_280 (
//    .x(16),
//    .d(u_2[279]),
//    .result(com_out[279])
//);

//compress_module compress_281 (
//    .x(16),
//    .d(u_2[280]),
//    .result(com_out[280])
//);

//compress_module compress_282 (
//    .x(16),
//    .d(u_2[281]),
//    .result(com_out[281])
//);

//compress_module compress_283 (
//    .x(16),
//    .d(u_2[282]),
//    .result(com_out[282])
//);

//compress_module compress_284 (
//    .x(16),
//    .d(u_2[283]),
//    .result(com_out[283])
//);

//compress_module compress_285 (
//    .x(16),
//    .d(u_2[284]),
//    .result(com_out[284])
//);

//compress_module compress_286 (
//    .x(16),
//    .d(u_2[285]),
//    .result(com_out[285])
//);

//compress_module compress_287 (
//    .x(16),
//    .d(u_2[286]),
//    .result(com_out[286])
//);

//compress_module compress_288 (
//    .x(16),
//    .d(u_2[287]),
//    .result(com_out[287])
//);

//compress_module compress_289 (
//    .x(16),
//    .d(u_2[288]),
//    .result(com_out[288])
//);

//compress_module compress_290 (
//    .x(16),
//    .d(u_2[289]),
//    .result(com_out[289])
//);

//compress_module compress_291 (
//    .x(16),
//    .d(u_2[290]),
//    .result(com_out[290])
//);

//compress_module compress_292 (
//    .x(16),
//    .d(u_2[291]),
//    .result(com_out[291])
//);

//compress_module compress_293 (
//    .x(16),
//    .d(u_2[292]),
//    .result(com_out[292])
//);

//compress_module compress_294 (
//    .x(16),
//    .d(u_2[293]),
//    .result(com_out[293])
//);

//compress_module compress_295 (
//    .x(16),
//    .d(u_2[294]),
//    .result(com_out[294])
//);

//compress_module compress_296 (
//    .x(16),
//    .d(u_2[295]),
//    .result(com_out[295])
//);

//compress_module compress_297 (
//    .x(16),
//    .d(u_2[296]),
//    .result(com_out[296])
//);

//compress_module compress_298 (
//    .x(16),
//    .d(u_2[297]),
//    .result(com_out[297])
//);

//compress_module compress_299 (
//    .x(16),
//    .d(u_2[298]),
//    .result(com_out[298])
//);

//compress_module compress_300 (
//    .x(16),
//    .d(u_2[299]),
//    .result(com_out[299])
//);

//compress_module compress_301 (
//    .x(16),
//    .d(u_2[300]),
//    .result(com_out[300])
//);

//compress_module compress_302 (
//    .x(16),
//    .d(u_2[301]),
//    .result(com_out[301])
//);

//compress_module compress_303 (
//    .x(16),
//    .d(u_2[302]),
//    .result(com_out[302])
//);

//compress_module compress_304 (
//    .x(16),
//    .d(u_2[303]),
//    .result(com_out[303])
//);

//compress_module compress_305 (
//    .x(16),
//    .d(u_2[304]),
//    .result(com_out[304])
//);

//compress_module compress_306 (
//    .x(16),
//    .d(u_2[305]),
//    .result(com_out[305])
//);

//compress_module compress_307 (
//    .x(16),
//    .d(u_2[306]),
//    .result(com_out[306])
//);

//compress_module compress_308 (
//    .x(16),
//    .d(u_2[307]),
//    .result(com_out[307])
//);

//compress_module compress_309 (
//    .x(16),
//    .d(u_2[308]),
//    .result(com_out[308])
//);

//compress_module compress_310 (
//    .x(16),
//    .d(u_2[309]),
//    .result(com_out[309])
//);

//compress_module compress_311 (
//    .x(16),
//    .d(u_2[310]),
//    .result(com_out[310])
//);

//compress_module compress_312 (
//    .x(16),
//    .d(u_2[311]),
//    .result(com_out[311])
//);

//compress_module compress_313 (
//    .x(16),
//    .d(u_2[312]),
//    .result(com_out[312])
//);

//compress_module compress_314 (
//    .x(16),
//    .d(u_2[313]),
//    .result(com_out[313])
//);

//compress_module compress_315 (
//    .x(16),
//    .d(u_2[314]),
//    .result(com_out[314])
//);

//compress_module compress_316 (
//    .x(16),
//    .d(u_2[315]),
//    .result(com_out[315])
//);

//compress_module compress_317 (
//    .x(16),
//    .d(u_2[316]),
//    .result(com_out[316])
//);

//compress_module compress_318 (
//    .x(16),
//    .d(u_2[317]),
//    .result(com_out[317])
//);

//compress_module compress_319 (
//    .x(16),
//    .d(u_2[318]),
//    .result(com_out[318])
//);

//compress_module compress_320 (
//    .x(16),
//    .d(u_2[319]),
//    .result(com_out[319])
//);

//compress_module compress_321 (
//    .x(16),
//    .d(u_2[320]),
//    .result(com_out[320])
//);

//compress_module compress_322 (
//    .x(16),
//    .d(u_2[321]),
//    .result(com_out[321])
//);

//compress_module compress_323 (
//    .x(16),
//    .d(u_2[322]),
//    .result(com_out[322])
//);

//compress_module compress_324 (
//    .x(16),
//    .d(u_2[323]),
//    .result(com_out[323])
//);

//compress_module compress_325 (
//    .x(16),
//    .d(u_2[324]),
//    .result(com_out[324])
//);

//compress_module compress_326 (
//    .x(16),
//    .d(u_2[325]),
//    .result(com_out[325])
//);

//compress_module compress_327 (
//    .x(16),
//    .d(u_2[326]),
//    .result(com_out[326])
//);

//compress_module compress_328 (
//    .x(16),
//    .d(u_2[327]),
//    .result(com_out[327])
//);

//compress_module compress_329 (
//    .x(16),
//    .d(u_2[328]),
//    .result(com_out[328])
//);

//compress_module compress_330 (
//    .x(16),
//    .d(u_2[329]),
//    .result(com_out[329])
//);

//compress_module compress_331 (
//    .x(16),
//    .d(u_2[330]),
//    .result(com_out[330])
//);

//compress_module compress_332 (
//    .x(16),
//    .d(u_2[331]),
//    .result(com_out[331])
//);

//compress_module compress_333 (
//    .x(16),
//    .d(u_2[332]),
//    .result(com_out[332])
//);

//compress_module compress_334 (
//    .x(16),
//    .d(u_2[333]),
//    .result(com_out[333])
//);

//compress_module compress_335 (
//    .x(16),
//    .d(u_2[334]),
//    .result(com_out[334])
//);

//compress_module compress_336 (
//    .x(16),
//    .d(u_2[335]),
//    .result(com_out[335])
//);

//compress_module compress_337 (
//    .x(16),
//    .d(u_2[336]),
//    .result(com_out[336])
//);

//compress_module compress_338 (
//    .x(16),
//    .d(u_2[337]),
//    .result(com_out[337])
//);

//compress_module compress_339 (
//    .x(16),
//    .d(u_2[338]),
//    .result(com_out[338])
//);

//compress_module compress_340 (
//    .x(16),
//    .d(u_2[339]),
//    .result(com_out[339])
//);

//compress_module compress_341 (
//    .x(16),
//    .d(u_2[340]),
//    .result(com_out[340])
//);

//compress_module compress_342 (
//    .x(16),
//    .d(u_2[341]),
//    .result(com_out[341])
//);

//compress_module compress_343 (
//    .x(16),
//    .d(u_2[342]),
//    .result(com_out[342])
//);

//compress_module compress_344 (
//    .x(16),
//    .d(u_2[343]),
//    .result(com_out[343])
//);

//compress_module compress_345 (
//    .x(16),
//    .d(u_2[344]),
//    .result(com_out[344])
//);

//compress_module compress_346 (
//    .x(16),
//    .d(u_2[345]),
//    .result(com_out[345])
//);

//compress_module compress_347 (
//    .x(16),
//    .d(u_2[346]),
//    .result(com_out[346])
//);

//compress_module compress_348 (
//    .x(16),
//    .d(u_2[347]),
//    .result(com_out[347])
//);

//compress_module compress_349 (
//    .x(16),
//    .d(u_2[348]),
//    .result(com_out[348])
//);

//compress_module compress_350 (
//    .x(16),
//    .d(u_2[349]),
//    .result(com_out[349])
//);

//compress_module compress_351 (
//    .x(16),
//    .d(u_2[350]),
//    .result(com_out[350])
//);

//compress_module compress_352 (
//    .x(16),
//    .d(u_2[351]),
//    .result(com_out[351])
//);

//compress_module compress_353 (
//    .x(16),
//    .d(u_2[352]),
//    .result(com_out[352])
//);

//compress_module compress_354 (
//    .x(16),
//    .d(u_2[353]),
//    .result(com_out[353])
//);

//compress_module compress_355 (
//    .x(16),
//    .d(u_2[354]),
//    .result(com_out[354])
//);

//compress_module compress_356 (
//    .x(16),
//    .d(u_2[355]),
//    .result(com_out[355])
//);

//compress_module compress_357 (
//    .x(16),
//    .d(u_2[356]),
//    .result(com_out[356])
//);

//compress_module compress_358 (
//    .x(16),
//    .d(u_2[357]),
//    .result(com_out[357])
//);

//compress_module compress_359 (
//    .x(16),
//    .d(u_2[358]),
//    .result(com_out[358])
//);

//compress_module compress_360 (
//    .x(16),
//    .d(u_2[359]),
//    .result(com_out[359])
//);

//compress_module compress_361 (
//    .x(16),
//    .d(u_2[360]),
//    .result(com_out[360])
//);

//compress_module compress_362 (
//    .x(16),
//    .d(u_2[361]),
//    .result(com_out[361])
//);

//compress_module compress_363 (
//    .x(16),
//    .d(u_2[362]),
//    .result(com_out[362])
//);

//compress_module compress_364 (
//    .x(16),
//    .d(u_2[363]),
//    .result(com_out[363])
//);

//compress_module compress_365 (
//    .x(16),
//    .d(u_2[364]),
//    .result(com_out[364])
//);

//compress_module compress_366 (
//    .x(16),
//    .d(u_2[365]),
//    .result(com_out[365])
//);

//compress_module compress_367 (
//    .x(16),
//    .d(u_2[366]),
//    .result(com_out[366])
//);

//compress_module compress_368 (
//    .x(16),
//    .d(u_2[367]),
//    .result(com_out[367])
//);

//compress_module compress_369 (
//    .x(16),
//    .d(u_2[368]),
//    .result(com_out[368])
//);

//compress_module compress_370 (
//    .x(16),
//    .d(u_2[369]),
//    .result(com_out[369])
//);

//compress_module compress_371 (
//    .x(16),
//    .d(u_2[370]),
//    .result(com_out[370])
//);

//compress_module compress_372 (
//    .x(16),
//    .d(u_2[371]),
//    .result(com_out[371])
//);

//compress_module compress_373 (
//    .x(16),
//    .d(u_2[372]),
//    .result(com_out[372])
//);

//compress_module compress_374 (
//    .x(16),
//    .d(u_2[373]),
//    .result(com_out[373])
//);

//compress_module compress_375 (
//    .x(16),
//    .d(u_2[374]),
//    .result(com_out[374])
//);

//compress_module compress_376 (
//    .x(16),
//    .d(u_2[375]),
//    .result(com_out[375])
//);

//compress_module compress_377 (
//    .x(16),
//    .d(u_2[376]),
//    .result(com_out[376])
//);

//compress_module compress_378 (
//    .x(16),
//    .d(u_2[377]),
//    .result(com_out[377])
//);

//compress_module compress_379 (
//    .x(16),
//    .d(u_2[378]),
//    .result(com_out[378])
//);

//compress_module compress_380 (
//    .x(16),
//    .d(u_2[379]),
//    .result(com_out[379])
//);

//compress_module compress_381 (
//    .x(16),
//    .d(u_2[380]),
//    .result(com_out[380])
//);

//compress_module compress_382 (
//    .x(16),
//    .d(u_2[381]),
//    .result(com_out[381])
//);

//compress_module compress_383 (
//    .x(16),
//    .d(u_2[382]),
//    .result(com_out[382])
//);

//compress_module compress_384 (
//    .x(16),
//    .d(u_2[383]),
//    .result(com_out[383])
//);

//compress_module compress_385 (
//    .x(16),
//    .d(u_2[384]),
//    .result(com_out[384])
//);

//compress_module compress_386 (
//    .x(16),
//    .d(u_2[385]),
//    .result(com_out[385])
//);

//compress_module compress_387 (
//    .x(16),
//    .d(u_2[386]),
//    .result(com_out[386])
//);

//compress_module compress_388 (
//    .x(16),
//    .d(u_2[387]),
//    .result(com_out[387])
//);

//compress_module compress_389 (
//    .x(16),
//    .d(u_2[388]),
//    .result(com_out[388])
//);

//compress_module compress_390 (
//    .x(16),
//    .d(u_2[389]),
//    .result(com_out[389])
//);

//compress_module compress_391 (
//    .x(16),
//    .d(u_2[390]),
//    .result(com_out[390])
//);

//compress_module compress_392 (
//    .x(16),
//    .d(u_2[391]),
//    .result(com_out[391])
//);

//compress_module compress_393 (
//    .x(16),
//    .d(u_2[392]),
//    .result(com_out[392])
//);

//compress_module compress_394 (
//    .x(16),
//    .d(u_2[393]),
//    .result(com_out[393])
//);

//compress_module compress_395 (
//    .x(16),
//    .d(u_2[394]),
//    .result(com_out[394])
//);

//compress_module compress_396 (
//    .x(16),
//    .d(u_2[395]),
//    .result(com_out[395])
//);

//compress_module compress_397 (
//    .x(16),
//    .d(u_2[396]),
//    .result(com_out[396])
//);

//compress_module compress_398 (
//    .x(16),
//    .d(u_2[397]),
//    .result(com_out[397])
//);

//compress_module compress_399 (
//    .x(16),
//    .d(u_2[398]),
//    .result(com_out[398])
//);

//compress_module compress_400 (
//    .x(16),
//    .d(u_2[399]),
//    .result(com_out[399])
//);

//compress_module compress_401 (
//    .x(16),
//    .d(u_2[400]),
//    .result(com_out[400])
//);

//compress_module compress_402 (
//    .x(16),
//    .d(u_2[401]),
//    .result(com_out[401])
//);

//compress_module compress_403 (
//    .x(16),
//    .d(u_2[402]),
//    .result(com_out[402])
//);

//compress_module compress_404 (
//    .x(16),
//    .d(u_2[403]),
//    .result(com_out[403])
//);

//compress_module compress_405 (
//    .x(16),
//    .d(u_2[404]),
//    .result(com_out[404])
//);

//compress_module compress_406 (
//    .x(16),
//    .d(u_2[405]),
//    .result(com_out[405])
//);

//compress_module compress_407 (
//    .x(16),
//    .d(u_2[406]),
//    .result(com_out[406])
//);

//compress_module compress_408 (
//    .x(16),
//    .d(u_2[407]),
//    .result(com_out[407])
//);

//compress_module compress_409 (
//    .x(16),
//    .d(u_2[408]),
//    .result(com_out[408])
//);

//compress_module compress_410 (
//    .x(16),
//    .d(u_2[409]),
//    .result(com_out[409])
//);

//compress_module compress_411 (
//    .x(16),
//    .d(u_2[410]),
//    .result(com_out[410])
//);

//compress_module compress_412 (
//    .x(16),
//    .d(u_2[411]),
//    .result(com_out[411])
//);

//compress_module compress_413 (
//    .x(16),
//    .d(u_2[412]),
//    .result(com_out[412])
//);

//compress_module compress_414 (
//    .x(16),
//    .d(u_2[413]),
//    .result(com_out[413])
//);

//compress_module compress_415 (
//    .x(16),
//    .d(u_2[414]),
//    .result(com_out[414])
//);

//compress_module compress_416 (
//    .x(16),
//    .d(u_2[415]),
//    .result(com_out[415])
//);

//compress_module compress_417 (
//    .x(16),
//    .d(u_2[416]),
//    .result(com_out[416])
//);

//compress_module compress_418 (
//    .x(16),
//    .d(u_2[417]),
//    .result(com_out[417])
//);

//compress_module compress_419 (
//    .x(16),
//    .d(u_2[418]),
//    .result(com_out[418])
//);

//compress_module compress_420 (
//    .x(16),
//    .d(u_2[419]),
//    .result(com_out[419])
//);

//compress_module compress_421 (
//    .x(16),
//    .d(u_2[420]),
//    .result(com_out[420])
//);

//compress_module compress_422 (
//    .x(16),
//    .d(u_2[421]),
//    .result(com_out[421])
//);

//compress_module compress_423 (
//    .x(16),
//    .d(u_2[422]),
//    .result(com_out[422])
//);

//compress_module compress_424 (
//    .x(16),
//    .d(u_2[423]),
//    .result(com_out[423])
//);

//compress_module compress_425 (
//    .x(16),
//    .d(u_2[424]),
//    .result(com_out[424])
//);

//compress_module compress_426 (
//    .x(16),
//    .d(u_2[425]),
//    .result(com_out[425])
//);

//compress_module compress_427 (
//    .x(16),
//    .d(u_2[426]),
//    .result(com_out[426])
//);

//compress_module compress_428 (
//    .x(16),
//    .d(u_2[427]),
//    .result(com_out[427])
//);

//compress_module compress_429 (
//    .x(16),
//    .d(u_2[428]),
//    .result(com_out[428])
//);

//compress_module compress_430 (
//    .x(16),
//    .d(u_2[429]),
//    .result(com_out[429])
//);

//compress_module compress_431 (
//    .x(16),
//    .d(u_2[430]),
//    .result(com_out[430])
//);

//compress_module compress_432 (
//    .x(16),
//    .d(u_2[431]),
//    .result(com_out[431])
//);

//compress_module compress_433 (
//    .x(16),
//    .d(u_2[432]),
//    .result(com_out[432])
//);

//compress_module compress_434 (
//    .x(16),
//    .d(u_2[433]),
//    .result(com_out[433])
//);

//compress_module compress_435 (
//    .x(16),
//    .d(u_2[434]),
//    .result(com_out[434])
//);

//compress_module compress_436 (
//    .x(16),
//    .d(u_2[435]),
//    .result(com_out[435])
//);

//compress_module compress_437 (
//    .x(16),
//    .d(u_2[436]),
//    .result(com_out[436])
//);

//compress_module compress_438 (
//    .x(16),
//    .d(u_2[437]),
//    .result(com_out[437])
//);

//compress_module compress_439 (
//    .x(16),
//    .d(u_2[438]),
//    .result(com_out[438])
//);

//compress_module compress_440 (
//    .x(16),
//    .d(u_2[439]),
//    .result(com_out[439])
//);

//compress_module compress_441 (
//    .x(16),
//    .d(u_2[440]),
//    .result(com_out[440])
//);

//compress_module compress_442 (
//    .x(16),
//    .d(u_2[441]),
//    .result(com_out[441])
//);

//compress_module compress_443 (
//    .x(16),
//    .d(u_2[442]),
//    .result(com_out[442])
//);

//compress_module compress_444 (
//    .x(16),
//    .d(u_2[443]),
//    .result(com_out[443])
//);

//compress_module compress_445 (
//    .x(16),
//    .d(u_2[444]),
//    .result(com_out[444])
//);

//compress_module compress_446 (
//    .x(16),
//    .d(u_2[445]),
//    .result(com_out[445])
//);

//compress_module compress_447 (
//    .x(16),
//    .d(u_2[446]),
//    .result(com_out[446])
//);

//compress_module compress_448 (
//    .x(16),
//    .d(u_2[447]),
//    .result(com_out[447])
//);

//compress_module compress_449 (
//    .x(16),
//    .d(u_2[448]),
//    .result(com_out[448])
//);

//compress_module compress_450 (
//    .x(16),
//    .d(u_2[449]),
//    .result(com_out[449])
//);

//compress_module compress_451 (
//    .x(16),
//    .d(u_2[450]),
//    .result(com_out[450])
//);

//compress_module compress_452 (
//    .x(16),
//    .d(u_2[451]),
//    .result(com_out[451])
//);

//compress_module compress_453 (
//    .x(16),
//    .d(u_2[452]),
//    .result(com_out[452])
//);

//compress_module compress_454 (
//    .x(16),
//    .d(u_2[453]),
//    .result(com_out[453])
//);

//compress_module compress_455 (
//    .x(16),
//    .d(u_2[454]),
//    .result(com_out[454])
//);

//compress_module compress_456 (
//    .x(16),
//    .d(u_2[455]),
//    .result(com_out[455])
//);

//compress_module compress_457 (
//    .x(16),
//    .d(u_2[456]),
//    .result(com_out[456])
//);

//compress_module compress_458 (
//    .x(16),
//    .d(u_2[457]),
//    .result(com_out[457])
//);

//compress_module compress_459 (
//    .x(16),
//    .d(u_2[458]),
//    .result(com_out[458])
//);

//compress_module compress_460 (
//    .x(16),
//    .d(u_2[459]),
//    .result(com_out[459])
//);

//compress_module compress_461 (
//    .x(16),
//    .d(u_2[460]),
//    .result(com_out[460])
//);

//compress_module compress_462 (
//    .x(16),
//    .d(u_2[461]),
//    .result(com_out[461])
//);

//compress_module compress_463 (
//    .x(16),
//    .d(u_2[462]),
//    .result(com_out[462])
//);

//compress_module compress_464 (
//    .x(16),
//    .d(u_2[463]),
//    .result(com_out[463])
//);

//compress_module compress_465 (
//    .x(16),
//    .d(u_2[464]),
//    .result(com_out[464])
//);

//compress_module compress_466 (
//    .x(16),
//    .d(u_2[465]),
//    .result(com_out[465])
//);

//compress_module compress_467 (
//    .x(16),
//    .d(u_2[466]),
//    .result(com_out[466])
//);

//compress_module compress_468 (
//    .x(16),
//    .d(u_2[467]),
//    .result(com_out[467])
//);

//compress_module compress_469 (
//    .x(16),
//    .d(u_2[468]),
//    .result(com_out[468])
//);

//compress_module compress_470 (
//    .x(16),
//    .d(u_2[469]),
//    .result(com_out[469])
//);

//compress_module compress_471 (
//    .x(16),
//    .d(u_2[470]),
//    .result(com_out[470])
//);

//compress_module compress_472 (
//    .x(16),
//    .d(u_2[471]),
//    .result(com_out[471])
//);

//compress_module compress_473 (
//    .x(16),
//    .d(u_2[472]),
//    .result(com_out[472])
//);

//compress_module compress_474 (
//    .x(16),
//    .d(u_2[473]),
//    .result(com_out[473])
//);

//compress_module compress_475 (
//    .x(16),
//    .d(u_2[474]),
//    .result(com_out[474])
//);

//compress_module compress_476 (
//    .x(16),
//    .d(u_2[475]),
//    .result(com_out[475])
//);

//compress_module compress_477 (
//    .x(16),
//    .d(u_2[476]),
//    .result(com_out[476])
//);

//compress_module compress_478 (
//    .x(16),
//    .d(u_2[477]),
//    .result(com_out[477])
//);

//compress_module compress_479 (
//    .x(16),
//    .d(u_2[478]),
//    .result(com_out[478])
//);

//compress_module compress_480 (
//    .x(16),
//    .d(u_2[479]),
//    .result(com_out[479])
//);

//compress_module compress_481 (
//    .x(16),
//    .d(u_2[480]),
//    .result(com_out[480])
//);

//compress_module compress_482 (
//    .x(16),
//    .d(u_2[481]),
//    .result(com_out[481])
//);

//compress_module compress_483 (
//    .x(16),
//    .d(u_2[482]),
//    .result(com_out[482])
//);

//compress_module compress_484 (
//    .x(16),
//    .d(u_2[483]),
//    .result(com_out[483])
//);

//compress_module compress_485 (
//    .x(16),
//    .d(u_2[484]),
//    .result(com_out[484])
//);

//compress_module compress_486 (
//    .x(16),
//    .d(u_2[485]),
//    .result(com_out[485])
//);

//compress_module compress_487 (
//    .x(16),
//    .d(u_2[486]),
//    .result(com_out[486])
//);

//compress_module compress_488 (
//    .x(16),
//    .d(u_2[487]),
//    .result(com_out[487])
//);

//compress_module compress_489 (
//    .x(16),
//    .d(u_2[488]),
//    .result(com_out[488])
//);

//compress_module compress_490 (
//    .x(16),
//    .d(u_2[489]),
//    .result(com_out[489])
//);

//compress_module compress_491 (
//    .x(16),
//    .d(u_2[490]),
//    .result(com_out[490])
//);

//compress_module compress_492 (
//    .x(16),
//    .d(u_2[491]),
//    .result(com_out[491])
//);

//compress_module compress_493 (
//    .x(16),
//    .d(u_2[492]),
//    .result(com_out[492])
//);

//compress_module compress_494 (
//    .x(16),
//    .d(u_2[493]),
//    .result(com_out[493])
//);

//compress_module compress_495 (
//    .x(16),
//    .d(u_2[494]),
//    .result(com_out[494])
//);

//compress_module compress_496 (
//    .x(16),
//    .d(u_2[495]),
//    .result(com_out[495])
//);

//compress_module compress_497 (
//    .x(16),
//    .d(u_2[496]),
//    .result(com_out[496])
//);

//compress_module compress_498 (
//    .x(16),
//    .d(u_2[497]),
//    .result(com_out[497])
//);

//compress_module compress_499 (
//    .x(16),
//    .d(u_2[498]),
//    .result(com_out[498])
//);

//compress_module compress_500 (
//    .x(16),
//    .d(u_2[499]),
//    .result(com_out[499])
//);

//compress_module compress_501 (
//    .x(16),
//    .d(u_2[500]),
//    .result(com_out[500])
//);

//compress_module compress_502 (
//    .x(16),
//    .d(u_2[501]),
//    .result(com_out[501])
//);

//compress_module compress_503 (
//    .x(16),
//    .d(u_2[502]),
//    .result(com_out[502])
//);

//compress_module compress_504 (
//    .x(16),
//    .d(u_2[503]),
//    .result(com_out[503])
//);

//compress_module compress_505 (
//    .x(16),
//    .d(u_2[504]),
//    .result(com_out[504])
//);

//compress_module compress_506 (
//    .x(16),
//    .d(u_2[505]),
//    .result(com_out[505])
//);

//compress_module compress_507 (
//    .x(16),
//    .d(u_2[506]),
//    .result(com_out[506])
//);

//compress_module compress_508 (
//    .x(16),
// +   .d(u_2[507]),
//    .result(com_out[507])
//);

//compress_module compress_509 (
//    .x(16),
//    .d(u_2[508]),
//    .result(com_out[508])
//);

//compress_module compress_510 (
//    .x(16),
//    .d(u_2[509]),
//    .result(com_out[509])
//);

//compress_module compress_511 (
//    .x(16),
//    .d(u_2[510]),
//    .result(com_out[510])
//);

//compress_module compress_512 (
//    .x(16),
//    .d(u_2[511]),
//    .result(com_out[511])
//);

         endmodule