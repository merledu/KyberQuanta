`timescale 1ns / 1ps
module encryption #( 
    parameter k = 3,
    parameter ELL = 16,
    parameter NUM_COEFFS = 256,
    parameter Q = 3329
)(
  input logic clk,
  input logic rst,
  input logic [7:0] pk[1183:0],    
  input logic [7:0] mess [32-1:0], 
  input [255:0] r,     
  output logic [15:0] A [0:2][0:2][0:255],
  output logic [ 16-1:0] T_hat_0 [0:256-1],
  output logic [ 16-1:0] T_hat_1 [0:256-1],
  output logic [ 16-1:0] T_hat_2 [0:256-1],
  output logic [ 16-1:0] m_dec [0:256-1],
  output logic [255:0] rho_t,
  output logic [11:0] y [0:2][255:0],
  output logic [11:0] e1 [0:2][255:0],
  output logic [11:0] e2 [255:0],
  output logic [15:0] y_ntt [0:2][255:0],
  output logic start_ntt,
  output logic start_inverse,
  output logic [15:0] mult_out_00 [255:0],
  output logic [15:0] mult_out_01 [255:0],
  output logic [15:0] mult_out_02 [255:0],
  output logic [15:0] mult_out_10 [255:0],
  output logic [15:0] mult_out_11 [255:0],
  output logic [15:0] mult_out_12 [255:0],
  output logic [15:0] mult_out_20 [255:0],
  output logic [15:0] mult_out_21 [255:0],
      output logic [15:0] mult_out_22 [255:0],
      output logic  done9_mul,
      output logic  done10_mul,
      output logic  done11_mul,
      output logic [15:0] mult_out_1 [255:0],
      output logic [15:0] mult_out_2 [255:0],
      output logic [15:0] mult_out_3 [255:0],
       output logic done0_mul,
        output logic  done1_mul,
       output  logic  done2_mul,
       output  logic  done3_mul,
       output  logic  done4_mul,
       output  logic  done5_mul,
       output  logic  done6_mul,
        output logic done7_mul,
        output logic  done8_mul,
        output logic start_mul, 
        output logic [15:0] mul_add [0:2][255:0],
        output logic [15:0] mul_add_t[0:2][255:0],           
         output   logic  done0_ntt,
          output  logic done1_ntt,
         output   logic done2_ntt,
            output logic done10_ntt,
               output logic done11_ntt,
               output logic done12_ntt,
               output logic [31:0] in_1 [256-1:0],
                 output logic [31:0] in_2 [256-1:0],
                 output logic [31:0] in_3 [256-1:0],
                 output logic [31:0] in_4 [256-1:0],
               output logic [31:0] in_5 [256-1:0],
           output logic [31:0] in_6 [256-1:0],
            output logic done13_ntt,
           output logic done14_ntt,
            output logic done15_ntt,
                 output logic [31:0] u [0:2][255:0] ,
                 output logic  [15:0] decom_out [0:256-1],
                 output logic [15:0] result [0:2][255:0],
                 output logic [15:0] com_out [0:2][255:0],
                 output logic [15:0] comp_v [0:2][255:0], 
                 output logic [7:0] encode_u [0:2] [320-1:0],
                 output logic [7:0] encode_v [0:2] [320-1:0]

      );
    

    logic [7:0] pk_slice0 [0:383];
    logic [7:0] pk_slice1 [0:383];
    logic [7:0] pk_slice2 [0:383];
    logic  done9_shake, done10_shake, done11_shake, done12_shake, done13_shake, done14_shake,done15_shake;
    logic  done0_cbd, done1_cbd, done2_cbd, done3_cbd, done4_cbd, done5_cbd,done6_cbd;
    logic [7:0] parse_array1 [767:0];
    logic [7:0] parse_array2 [767:0];
    logic [7:0] parse_array3 [767:0];
    logic [7:0] parse_array4 [767:0];
    logic [7:0] parse_array5 [767:0];
    logic [7:0] parse_array6 [767:0];
    logic [7:0] parse_array7 [767:0];
    logic [7:0] parse_array8 [767:0];
    logic [7:0] parse_array9 [767:0];
    logic start1;
    logic done0, done1, done2, done3, done4, done5, done6, done7, done8, done9;
    logic done0_shake,done1_shake,done2_shake,done3_shake,done4_shake,done5_shake,done6_shake,done7_shake,done8_shake;
    logic all_shake_done;
    logic [7:0] prf_bytes_0 [127:0];
    logic [7:0] prf_bytes_1 [127:0];
    logic [7:0] prf_bytes_2 [127:0];
    logic [7:0] prf_bytes_3 [127:0];
    logic [7:0] prf_bytes_4 [127:0];
    logic [7:0] prf_bytes_5 [127:0];
    logic [7:0] prf_bytes_6 [127:0];
    logic [1023:0] prf_0, prf_1, prf_2, prf_3, prf_4, prf_5, prf_6;
    logic  start_parse, start_cbd, start_prf;
    logic [15:0] zetas [127:0];
    logic ntt_started;
    logic mul;
    logic [268-1:0] r0;
    logic [268-1:0] r1;
    logic [268-1:0] r2;
    logic [268-1:0] r3;
    logic [268-1:0] r4;
    logic [268-1:0] r5;
   

    
    
    assign pk_slice0 = pk[383:0];
    assign pk_slice1 = pk[767:384];
    assign pk_slice2 = pk[1151:768];
   
assign rho_t = {
           pk[1152], pk[1153], pk[1154], pk[1155],
           pk[1156], pk[1157], pk[1158], pk[1159],
           pk[1160], pk[1161], pk[1162], pk[1163],
           pk[1164], pk[1165], pk[1166], pk[1167],
           pk[1168], pk[1169], pk[1170], pk[1171],
           pk[1172], pk[1173], pk[1174], pk[1175],
           pk[1176], pk[1177], pk[1178], pk[1179],
           pk[1180], pk[1181], pk[1182], pk[1183]
       };


    decode #(.ELL(16), .NUM_COEFFS(256), .BYTE_COUNT(384)) dec0 (
        .byte_array(pk_slice0),
        .len(384),
        .coeffs(T_hat_0)
    );

    decode #(.ELL(16), .NUM_COEFFS(256), .BYTE_COUNT(384)) dec1 (
        .byte_array(pk_slice1),
        .len(384),
        .coeffs(T_hat_1)
    );

    decode #(.ELL(16), .NUM_COEFFS(256), .BYTE_COUNT(384)) dec2 (
        .byte_array(pk_slice2),
        .len(384),
        .coeffs(T_hat_2)
    );
   logic [7:0] mess [32-1:0];
    assign mess[0]  = 8'hEB;
   assign mess[1]  = 8'h4A;
   assign mess[2]  = 8'h7C;
   assign mess[3]  = 8'h66;
   assign mess[4]  = 8'hEF;
   assign mess[5]  = 8'h4E;
   assign mess[6]  = 8'hBA;
   assign mess[7]  = 8'h2D;
   assign mess[8]  = 8'hDB;
   assign mess[9]  = 8'h38;
   assign mess[10] = 8'hC8;
   assign mess[11] = 8'h8D;
   assign mess[12] = 8'h8B;
   assign mess[13] = 8'hC7;
   assign mess[14] = 8'h06;
   assign mess[15] = 8'hB1;
   assign mess[16] = 8'hD6;
   assign mess[17] = 8'h39;
   assign mess[18] = 8'h00;
   assign mess[19] = 8'h21;
   assign mess[20] = 8'h98;
   assign mess[21] = 8'h17;
   assign mess[22] = 8'h2A;
   assign mess[23] = 8'h7B;
   assign mess[24] = 8'h19;
   assign mess[25] = 8'h42;
   assign mess[26] = 8'hEC;
   assign mess[27] = 8'hA8;
   assign mess[28] = 8'hF6;
   assign mess[29] = 8'hC0;
   assign mess[30] = 8'h01;
   assign mess[31] = 8'hBA;

  decode #(.ELL(16), .NUM_COEFFS(256),.BYTE_COUNT(32)) dec4 (
                         .byte_array(mess),
                         .len(32),
                         .coeffs(m_dec)
                     );     
              //--------------------------XOF 1--------------------------------------
    logic [276-1:0] datain;
    logic [6144-1:0] xof;
    
   assign datain = {4'hF,8'h00, 8'h00,rho_t};
   assign message = datain; 
//   assign done0_shake = 1'b1;
    sponge #(
     .msg_len(276),
     .d_len(6144),
     .capacity(256),
     .r(1600 - 256)
 ) shake1(
        .clk(clk),
        .reset(rst),
        .start(start1),
        .message(datain),
        .z(xof),
        .done(done0_shake)
    );
            
           
           //--------------------------XOF 2--------------------------------------
              logic [276-1:0] datain2;
                   logic [6144-1:0] xof2;
//                  assign message = datain2; 
                   assign datain2 = {4'hF ,8'h00, 8'h02,rho_t};     
                    
                   sponge #(
                    .msg_len(276),
                    .d_len(6144),
                    .capacity(256),
                    .r(1600 - 256)
                ) shake2(
                       .clk(clk),
                       .reset(rst),
                       .start(start1),
                       .message(datain2),
                       .z(xof2),
                       .done(done1_shake)
                   ); 
                    
                 //--------------------------XOF 3--------------------------------------
               logic [276-1:0] datain3;
               logic [6144-1:0] xof3;
//                        assign message = datain3;                           
               assign datain3 = {4'hF , 8'h00, 8'h11,rho_t };      
               sponge #(
                    .msg_len(276),
                     .d_len(6144),
                     .capacity(256),
                     .r(1600 - 256)
                                  ) shake3(
                                        .clk(clk),
                                         .reset(rst),
                                         .start(start1),
                                        .message(datain3),
                                          .z(xof3),
                                           .done(done2_shake)
                                                  );
   
                    // --------------------------XOF 4--------------------------------------
              logic [276-1:0] datain4;
              logic [6144-1:0] xof4;
//                                                            assign message = datain4; 
              assign datain4 = {4'hF ,  8'h01 , 8'h00,rho_t };
              sponge #(
                        .msg_len(276),
                         .d_len(6144),
                         .capacity(256),
                         .r(1600 - 256)
                   ) shake4 (
                              .clk(clk),
                             .reset(rst),
                             .start(start1),
                            .message(datain4),
                             .z(xof4),
                             .done( done3_shake)
                                        );        
                  
                    // --------------------------XOF 5--------------------------------------
                         logic [276-1:0] datain5;
                  logic [6144-1:0] xof5;
//                assign message = datain5; 
            assign datain5 = {4'hF ,  8'h01 , 8'h01,rho_t };
        sponge #(
                      .msg_len(276),
                      .d_len(6144),
                      .capacity(256),
                       .r(1600 - 256)
                                       )
                 shake5 (
                         .clk(clk),
                         .reset(rst),
                         .start(start1),
                         .message(datain5),
                         .z(xof5),
                         .done( done4_shake)
                          );  
                 
                    // --------------------------XOF 6--------------------------------------
                       logic [276-1:0] datain6;
                       logic [6144-1:0] xof6;
//                       assign message = datain6; 
                       assign datain6 = {4'hF ,  8'h1 , 8'h2,rho_t };
                       sponge #(
                       .msg_len(276),
                       .d_len(6144),
                       .capacity(256),
                       .r(1600 - 256)
                       ) shake6 (
                       .clk(clk),
                        .reset(rst),
                        .start(start1),
                        .message(datain6),
                        .z(xof6),
                        .done( done5_shake)
                        );
                  
               // --------------------------XOF 7--------------------------------------
                   logic [276-1:0] datain7;
                   logic [6144-1:0] xof7;
//                    assign message = datain7; 
                   assign datain7 = {4'hF ,  8'h02 , 8'h00,rho_t };
                   sponge #(
                   .msg_len(276),
                   .d_len(6144),
                   .capacity(256),
                   .r(1600 - 256)
                   ) shake7 (
                   .clk(clk),
                   .reset(rst),
                   .start(start1),
                   .message(datain7),
                   .z(xof7),
                   .done( done6_shake)
                    );
   
                    // --------------------------XOF 8--------------------------------------
                     logic [276-1:0] datain8;
                     logic [6144-1:0] xof8;
//                     assign message = datain8; 
                     assign datain8 = {4'hF ,  8'h02 , 8'h01,rho_t };
                      sponge #(
                       .msg_len(276),
                       .d_len(6144),
                       .capacity(256),
                        .r(1600 - 256)
                         ) shake8 (
                          .clk(clk),
                           .reset(rst),
                            .start(start1),
                            .message(datain8),
                            .z(xof8),
                             .done( done7_shake)
                              );
                                                                                                          
                                                                                                          // --------------------------XOF 9--------------------------------------
          logic [276-1:0] datain9;
          logic [6144-1:0] xof9;
//        assign message = datain9; 
          assign datain9 = {4'hF ,  8'h2 , 8'h2,rho_t };
          sponge #(
           .msg_len(276),
           .d_len(6144),
           .capacity(256),
           .r(1600 - 256)
            ) shake9 (
            .clk(clk),
            .reset(rst),
            .start(start1),
            .message(datain9),
            .z(xof9),
            .done( done8_shake)
             );
       parse parse_00 (.clk(clk),.rst(rst),.start(done0_shake),.done(done0), .B(parse_array1), .a(A[0][0]));
       parse parse_01 (.clk(clk),.rst(rst),.start(done1_shake),.done(done1),.B(parse_array2), .a(A[0][1]));
       parse parse_02 (.clk(clk),.rst(rst),.start(done2_shake),.done(done2),.B(parse_array3), .a(A[0][2]));
       
       parse parse_10 (.clk(clk),.rst(rst),.start(done3_shake),.done(done3),.B(parse_array4), .a(A[1][0]));
       parse parse_11 (.clk(clk),.rst(rst),.start(done4_shake),.done(done4),.B(parse_array5), .a(A[1][1]));
       parse parse_12 (.clk(clk),.rst(rst),.start(done4_shake),.done(done5),.B(parse_array6), .a(A[1][2]));
       
       parse parse_20 (.clk(clk),.rst(rst),.start(done4_shake),.done(done6),.B(parse_array7), .a(A[2][0]));
       parse parse_21 (.clk(clk),.rst(rst),.start(done4_shake),.done(done7),.B(parse_array8), .a(A[2][1]));
       parse parse_22 (.clk(clk),.rst(rst),.start(done8_shake),.done(done8),.B(parse_array9), .a(A[2][2]));
       

     
//     //-----------------prf0-------------------------
    
     
     assign r0 = {4'h1111, 8'h00,r}; 
     assign r1 = {4'h1111, 8'h01,r};
      assign r2 = {4'h1111, 8'h02,r};
         assign r3 = {4'h1111, 8'h03,r};  
            assign r4 = {4'h1111, 8'h04,r}; 
             assign r5 = {4'h1111, 8'h05,r};
             
     sponge #(.msg_len(268),
      .d_len(1024), 
      .capacity(512),
       .r(1600 - 512))
        prf0 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r0),
         .z(prf_0),
         .done(done9_shake)
     );
     
  
     sponge #(.msg_len(268), 
     .d_len(1024), 
     .capacity(512), 
     .r(1600 - 512)) 
     prf1 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r1),
         .z(prf_1),
         .done(done10_shake)
     );
     
    
     sponge #(.msg_len(268), 
     .d_len(1024), 
     .capacity(512),
      .r(1600 - 512)) 
      prf2 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r2),
         .z(prf_2),
         .done(done11_shake)
     );
   
  
     sponge #(.msg_len(268),
      .d_len(1024), 
      .capacity(512),
       .r(1600 - 512))
        prf3 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r3),
         .z(prf_3),
         .done(done12_shake)
     );
     
   
     sponge #(.msg_len(268),
      .d_len(1024),
       .capacity(512),
        .r(1600 - 512)) 
        prf4 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r4),
         .z(prf_4),
         .done(done13_shake)
     );
     
     
    
     sponge #(.msg_len(268),
      .d_len(1024),
       .capacity(512),
        .r(1600 - 512))
      prf5 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r5),
         .z(prf_5),
         .done(done14_shake)
     );
                  
        CBD cbd0 (.clk(clk), .reset(rst), .start(done14_shake), .done(done0_cbd), .byte_array(prf_bytes_0), .len(128), .f(y[0]));
        CBD cbd1 (.clk(clk), .reset(rst), .start(done14_shake), .done(done1_cbd), .byte_array(prf_bytes_1), .len(128), .f(y[1]));
        CBD cbd2 (.clk(clk), .reset(rst), .start(done14_shake), .done(done2_cbd), .byte_array(prf_bytes_2), .len(128), .f(y[2]));
        
        CBD cbd3 (.clk(clk), .reset(rst), .start(done14_shake), .done(done3_cbd), .byte_array(prf_bytes_3), .len(128), .f(e1[0]));
        CBD cbd4 (.clk(clk), .reset(rst), .start(done14_shake), .done(done4_cbd), .byte_array(prf_bytes_4), .len(128), .f(e1[1]));
        CBD cbd5 (.clk(clk), .reset(rst), .start(done14_shake), .done(done5_cbd), .byte_array(prf_bytes_5), .len(128), .f(e1[2]));
        

        logic [268-1:0] r6;
        assign r6 = {4'h1111, 8'h06,r}; 
        sponge #(.msg_len(268),
             .d_len(1024), 
             .capacity(512),
              .r(1600 - 512))
               prf6 (
                .clk(clk),
                .reset(rst),
                .start(done8),
                .message(r6),
                .z(prf_6),
                .done(done15_shake)
            );
               CBD cbd6  (
                  .clk(clk), 
                           .reset(rst), 
                           .start(done14_shake), 
                           .done(done6_cbd), 
                           .byte_array(prf_bytes_6), 
                           .len(128), 
                           .f(e2)
              );
              
               assign start_ntt = (done5_cbd && !done0_ntt && !done1_ntt && !done2_ntt);
               
                   ntt ntt_y0 (.clk(clk), .reset(rst), .f(y[0]), .start(start_ntt), .done(done0_ntt), .f_hat(y_ntt[0]));
                   ntt ntt_y1 (.clk(clk), .reset(rst), .f(y[1]), .start(start_ntt), .done(done1_ntt),.f_hat(y_ntt[1]));
                   ntt ntt_y2 (.clk(clk), .reset(rst), .f(y[2]), .start(start_ntt), .done(done2_ntt),.f_hat(y_ntt[2]));
           
                      
                     assign start_mul = (done0_ntt && done1_ntt && done2_ntt);
                  
                      multiply_ntts mul_00 (.clk(clk), .reset(rst),.f(A[0][0]), .g(y_ntt[0]), .zetas(zetas), .h(mult_out_00), .start(start_mul), .done(done0_mul));
                      multiply_ntts mul_01 (.clk(clk), .reset(rst),.f(A[0][1]), .g(y_ntt[1]), .zetas(zetas), .h(mult_out_01),.start(start_mul), .done(done1_mul));
                      multiply_ntts mul_02 (.clk(clk), .reset(rst),.f(A[0][2]), .g(y_ntt[2]), .zetas(zetas), .h(mult_out_02),.start(start_mul), .done(done2_mul));
                  
                      multiply_ntts mul_10 (.clk(clk), .reset(rst),.f(A[1][0]), .g(y_ntt[0]), .zetas(zetas), .h(mult_out_10), .start(start_mul), .done(done3_mul));
                      multiply_ntts mul_11 (.clk(clk), .reset(rst),.f(A[1][1]), .g(y_ntt[1]),.zetas(zetas), .h(mult_out_11), .start(start_mul), .done(done4_mul));
                      multiply_ntts mul_12 (.clk(clk), .reset(rst),.f(A[1][2]), .g(y_ntt[2]), .zetas(zetas),.h(mult_out_12), .start(start_mul), .done(done5_mul));
                  
                      multiply_ntts mul_20 (.clk(clk), .reset(rst),.f(A[2][0]), .g(y_ntt[0]),.zetas(zetas), .h(mult_out_20), .start(start_mul),.done(done6_mul));
                      multiply_ntts mul_21 (.clk(clk), .reset(rst),.f(A[2][1]), .g(y_ntt[1]), .zetas(zetas),.h(mult_out_21), .start(start_mul), .done(done7_mul));
                      multiply_ntts mul_22 (.clk(clk), .reset(rst),.f(A[2][2]), .g(y_ntt[2]), .zetas(zetas),.h(mult_out_22), .start(start_mul), .done(done8_mul));

                      
                      multiply_ntts
                          mult_1 (
                              .clk(clk),
                              .reset(rst),
                              .f(T_hat_0),  // T_hat_0_16 is a 16-bit array
                              .g(y_ntt[0]),  // y_ntt_0_16 is now a 1D array
                              .zetas(zetas),
                              .h(mult_out_1),
                              .start(start_mul),
                              .done(done9_mul)
                          );
                      
                      multiply_ntts
                          mult_2 (
                              .clk(clk),
                              .reset(rst),
                              .f(T_hat_1),  // T_hat_1_16 is a 16-bit array
                              .g(y_ntt[1]),  // y_ntt_1_16 is now a 1D array
                              .zetas(zetas),
                              .h(mult_out_2),
                              .start(start_mul),
                              .done(done10_mul)
                          );
                      
                      multiply_ntts
                          mult_3 (
                              .clk(clk),
                              .reset(rst),
                              .f(T_hat_2),  
                              .g(y_ntt[2]),  
                              .zetas(zetas),
                              .h(mult_out_3),
                              .start(start_mul),
                              .done(done11_mul)
                          );
                          assign start_inverse = (done3_mul && done4_mul && done5_mul );
                          
                          ////AT x Y inverse
//                          logic  [31:0] in_1 [256-1:0];
                          
                          inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_1 (
                              .clk(clk),
                              .rst(rst),
                              .f(mul_add[0]),
                              .start_ntt(start_inverse),
                              .done_ntt(done10_ntt),
                              .f_hat(in_1)
                          );
                          
                          inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_2 (
                              .clk(clk),
                              .rst(rst),
                              .f(mul_add[1]),
                              .start_ntt(start_inverse),
                              .done_ntt(done11_ntt),
                              .f_hat(in_2)
                          );
                          
                          inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_3 (
                              .clk(clk),
                              .rst(rst),
                              .f(mul_add[2]),
                              .start_ntt(start_inverse),
                              .done_ntt(done12_ntt),
                              .f_hat(in_3)
                          );
                           inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_4 (
                                                       .clk(clk),
                                                       .rst(rst),
                                                       .f(mul_add_t[0]),
                                                       .start_ntt(start_inverse),
                                                       .done_ntt(done13_ntt),
                                                       .f_hat(in_4)
                                                   );
                                                   
                        inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_5 (
                                                       .clk(clk),
                                                       .rst(rst),
                                                       .f(mul_add_t[1]),
                                                       .start_ntt(start_inverse),
                                                       .done_ntt(done14_ntt),
                                                       .f_hat(in_5)
                                                   );
                                                   
                        inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_6 (
                                                       .clk(clk),
                                                       .rst(rst),
                                                       .f(mul_add_t[2]),
                                                       .start_ntt(start_inverse),
                                                       .done_ntt(done15_ntt),
                                                       .f_hat(in_6)
                                                   );
                           

                      decompress_module decompress_inst0 (
                                            .x(m_dec[0]),
                                            .d(16),
                                            .result(decom_out[0])
                                        );
                                        
                                        decompress_module decompress_inst1 (
                                            .x(m_dec[1]),
                                            .d(16),
                                            .result(decom_out[1])
                                        );
                                        
                                        decompress_module decompress_inst2 (
                                            .x(m_dec[2]),
                                            .d(16),
                                            .result(decom_out[2])
                                        );
                                        
                                        decompress_module decompress_inst3 (
                                            .x(m_dec[3]),
                                            .d(16),
                                            .result(decom_out[3])
                                        );
                                        
                                        decompress_module decompress_inst4 (
                                            .x(m_dec[4]),
                                            .d(16),
                                            .result(decom_out[4])
                                        );
                                        
                                        decompress_module decompress_inst5 (
                                            .x(m_dec[5]),
                                            .d(16),
                                            .result(decom_out[5])
                                        );
                                        
                                        decompress_module decompress_inst6 (
                                            .x(m_dec[6]),
                                            .d(16),
                                            .result(decom_out[6])
                                        );
                                        
                                        decompress_module decompress_inst7 (
                                            .x(m_dec[7]),
                                            .d(16),
                                            .result(decom_out[7])
                                        );
                                        
                                        decompress_module decompress_inst8 (
                                            .x(m_dec[8]),
                                            .d(16),
                                            .result(decom_out[8])
                                        );
                                        
                                        decompress_module decompress_inst9 (
                                            .x(m_dec[9]),
                                            .d(16),
                                            .result(decom_out[9])
                                        );
                                        
                                        decompress_module decompress_inst10 (
                                            .x(m_dec[10]),
                                            .d(16),
                                            .result(decom_out[10])
                                        );
                                        
                                        decompress_module decompress_inst11 (
                                            .x(m_dec[11]),
                                            .d(16),
                                            .result(decom_out[11])
                                        );
                                        
                                        decompress_module decompress_inst12 (
                                            .x(m_dec[12]),
                                            .d(16),
                                            .result(decom_out[12])
                                        );
                                        
                                        decompress_module decompress_inst13 (
                                            .x(m_dec[13]),
                                            .d(16),
                                            .result(decom_out[13])
                                        );
                                        
                                        decompress_module decompress_inst14 (
                                            .x(m_dec[14]),
                                            .d(16),
                                            .result(decom_out[14])
                                        );
                                        
                                        decompress_module decompress_inst15 (
                                            .x(m_dec[15]),
                                            .d(16),
                                            .result(decom_out[15])
                                        );
                                        
                                        decompress_module decompress_inst16 (
                                            .x(m_dec[16]),
                                            .d(16),
                                            .result(decom_out[16])
                                        );
                                        
                                        decompress_module decompress_inst17 (
                                            .x(m_dec[17]),
                                            .d(16),
                                            .result(decom_out[17])
                                        );
                                        
                                        decompress_module decompress_inst18 (
                                            .x(m_dec[18]),
                                            .d(16),
                                            .result(decom_out[18])
                                        );
                                        
                                        decompress_module decompress_inst19 (
                                            .x(m_dec[19]),
                                            .d(16),
                                            .result(decom_out[19])
                                        );
                                        
                                        decompress_module decompress_inst20 (
                                            .x(m_dec[20]),
                                            .d(16),
                                            .result(decom_out[20])
                                        );
                                        
                                        decompress_module decompress_inst21 (
                                            .x(m_dec[21]),
                                            .d(16),
                                            .result(decom_out[21])
                                        );
                                        
                                        decompress_module decompress_inst22 (
                                            .x(m_dec[22]),
                                            .d(16),
                                            .result(decom_out[22])
                                        );
                                        
                                        decompress_module decompress_inst23 (
                                            .x(m_dec[23]),
                                            .d(16),
                                            .result(decom_out[23])
                                        );
                                        
                                        decompress_module decompress_inst24 (
                                            .x(m_dec[24]),
                                            .d(16),
                                            .result(decom_out[24])
                                        );
                                        
                                        decompress_module decompress_inst25 (
                                            .x(m_dec[25]),
                                            .d(16),
                                            .result(decom_out[25])
                                        );
                                        
                                        decompress_module decompress_inst26 (
                                            .x(m_dec[26]),
                                            .d(16),
                                            .result(decom_out[26])
                                        );
                                        
                                        decompress_module decompress_inst27 (
                                            .x(m_dec[27]),
                                            .d(16),
                                            .result(decom_out[27])
                                        );
                                        
                                        decompress_module decompress_inst28 (
                                            .x(m_dec[28]),
                                            .d(16),
                                            .result(decom_out[28])
                                        );
                                        
                                        decompress_module decompress_inst29 (
                                            .x(m_dec[29]),
                                            .d(16),
                                            .result(decom_out[29])
                                        );
                                        
                                        decompress_module decompress_inst30 (
                                            .x(m_dec[30]),
                                            .d(16),
                                            .result(decom_out[30])
                                        );
                                        
                                        decompress_module decompress_inst31 (
                                            .x(m_dec[31]),
                                            .d(16),
                                            .result(decom_out[31])
                                        );
                                        
                                        decompress_module decompress_inst32 (
                                            .x(m_dec[32]),
                                            .d(16),
                                            .result(decom_out[32])
                                        );
                                        
                                        decompress_module decompress_inst33 (
                                            .x(m_dec[33]),
                                            .d(16),
                                            .result(decom_out[33])
                                        );
                                        
                                        decompress_module decompress_inst34 (
                                            .x(m_dec[34]),
                                            .d(16),
                                            .result(decom_out[34])
                                        );
                                        
                                        decompress_module decompress_inst35 (
                                            .x(m_dec[35]),
                                            .d(16),
                                            .result(decom_out[35])
                                        );
                                        
                                        decompress_module decompress_inst36 (
                                            .x(m_dec[36]),
                                            .d(16),
                                            .result(decom_out[36])
                                        );
                                        
                                        decompress_module decompress_inst37 (
                                            .x(m_dec[37]),
                                            .d(16),
                                            .result(decom_out[37])
                                        );
                                        
                                        decompress_module decompress_inst38 (
                                            .x(m_dec[38]),
                                            .d(16),
                                            .result(decom_out[38])
                                        );
                                        
                                        decompress_module decompress_inst39 (
                                            .x(m_dec[39]),
                                            .d(16),
                                            .result(decom_out[39])
                                        );
                                        
                                        decompress_module decompress_inst40 (
                                            .x(m_dec[40]),
                                            .d(16),
                                            .result(decom_out[40])
                                        );
                                        
                                        decompress_module decompress_inst41 (
                                            .x(m_dec[41]),
                                            .d(16),
                                            .result(decom_out[41])
                                        );
                                        
                                        decompress_module decompress_inst42 (
                                            .x(m_dec[42]),
                                            .d(16),
                                            .result(decom_out[42])
                                        );
                                        
                                        decompress_module decompress_inst43 (
                                            .x(m_dec[43]),
                                            .d(16),
                                            .result(decom_out[43])
                                        );
                                        
                                        decompress_module decompress_inst44 (
                                            .x(m_dec[44]),
                                            .d(16),
                                            .result(decom_out[44])
                                        );
                                        
                                        decompress_module decompress_inst45 (
                                            .x(m_dec[45]),
                                            .d(16),
                                            .result(decom_out[45])
                                        );
                                        
                                        decompress_module decompress_inst46 (
                                            .x(m_dec[46]),
                                            .d(16),
                                            .result(decom_out[46])
                                        );
                                        
                                        decompress_module decompress_inst47 (
                                            .x(m_dec[47]),
                                            .d(16),
                                            .result(decom_out[47])
                                        );
                                        
                                        decompress_module decompress_inst48 (
                                            .x(m_dec[48]),
                                            .d(16),
                                            .result(decom_out[48])
                                        );
                                        
                                        decompress_module decompress_inst49 (
                                            .x(m_dec[49]),
                                            .d(16),
                                            .result(decom_out[49])
                                        );
                                        
                                        decompress_module decompress_inst50 (
                                            .x(m_dec[50]),
                                            .d(16),
                                            .result(decom_out[50])
                                        );
                                        
                                        decompress_module decompress_inst51 (
                                            .x(m_dec[51]),
                                            .d(16),
                                            .result(decom_out[51])
                                        );
                                        
                                        decompress_module decompress_inst52 (
                                            .x(m_dec[52]),
                                            .d(16),
                                            .result(decom_out[52])
                                        );
                                        
                                        decompress_module decompress_inst53 (
                                            .x(m_dec[53]),
                                            .d(16),
                                            .result(decom_out[53])
                                        );
                                        
                                        decompress_module decompress_inst54 (
                                            .x(m_dec[54]),
                                            .d(16),
                                            .result(decom_out[54])
                                        );
                                        
                                        decompress_module decompress_inst55 (
                                            .x(m_dec[55]),
                                            .d(16),
                                            .result(decom_out[55])
                                        );
                                        
                                        decompress_module decompress_inst56 (
                                            .x(m_dec[56]),
                                            .d(16),
                                            .result(decom_out[56])
                                        );
                                        
                                        decompress_module decompress_inst57 (
                                            .x(m_dec[57]),
                                            .d(16),
                                            .result(decom_out[57])
                                        );
                                        
                                        decompress_module decompress_inst58 (
                                            .x(m_dec[58]),
                                            .d(16),
                                            .result(decom_out[58])
                                        );
                                        
                                        decompress_module decompress_inst59 (
                                            .x(m_dec[59]),
                                            .d(16),
                                            .result(decom_out[59])
                                        );
                                        
                                        decompress_module decompress_inst60 (
                                            .x(m_dec[60]),
                                            .d(16),
                                            .result(decom_out[60])
                                        );
                                        
                                        decompress_module decompress_inst61 (
                                            .x(m_dec[61]),
                                            .d(16),
                                            .result(decom_out[61])
                                        );
                                        
                                        decompress_module decompress_inst62 (
                                            .x(m_dec[62]),
                                            .d(16),
                                            .result(decom_out[62])
                                        );
                                        
                                        decompress_module decompress_inst63 (
                                            .x(m_dec[63]),
                                            .d(16),
                                            .result(decom_out[63])
                                        );
                                        
                                        decompress_module decompress_inst64 (
                                            .x(m_dec[64]),
                                            .d(16),
                                            .result(decom_out[64])
                                        );
                                        
                                        decompress_module decompress_inst65 (
                                            .x(m_dec[65]),
                                            .d(16),
                                            .result(decom_out[65])
                                        );
                                        
                                        decompress_module decompress_inst66 (
                                            .x(m_dec[66]),
                                            .d(16),
                                            .result(decom_out[66])
                                        );
                                        
                                        decompress_module decompress_inst67 (
                                            .x(m_dec[67]),
                                            .d(16),
                                            .result(decom_out[67])
                                        );
                                        
                                        decompress_module decompress_inst68 (
                                            .x(m_dec[68]),
                                            .d(16),
                                            .result(decom_out[68])
                                        );
                                        
                                        decompress_module decompress_inst69 (
                                            .x(m_dec[69]),
                                            .d(16),
                                            .result(decom_out[69])
                                        );
                                        
                                        decompress_module decompress_inst70 (
                                            .x(m_dec[70]),
                                            .d(16),
                                            .result(decom_out[70])
                                        );
                                        
                                        decompress_module decompress_inst71 (
                                            .x(m_dec[71]),
                                            .d(16),
                                            .result(decom_out[71])
                                        );
                                        
                                        decompress_module decompress_inst72 (
                                            .x(m_dec[72]),
                                            .d(16),
                                            .result(decom_out[72])
                                        );
                                        
                                        decompress_module decompress_inst73 (
                                            .x(m_dec[73]),
                                            .d(16),
                                            .result(decom_out[73])
                                        );
                                        
                                        decompress_module decompress_inst74 (
                                            .x(m_dec[74]),
                                            .d(16),
                                            .result(decom_out[74])
                                        );
                                        
                                        decompress_module decompress_inst75 (
                                            .x(m_dec[75]),
                                            .d(16),
                                            .result(decom_out[75])
                                        );
                                        
                                        decompress_module decompress_inst76 (
                                            .x(m_dec[76]),
                                            .d(16),
                                            .result(decom_out[76])
                                        );
                                        
                                        decompress_module decompress_inst77 (
                                            .x(m_dec[77]),
                                            .d(16),
                                            .result(decom_out[77])
                                        );
                                        
                                        decompress_module decompress_inst78 (
                                            .x(m_dec[78]),
                                            .d(16),
                                            .result(decom_out[78])
                                        );
                                        
                                        decompress_module decompress_inst79 (
                                            .x(m_dec[79]),
                                            .d(16),
                                            .result(decom_out[79])
                                        );
                                        
                                        decompress_module decompress_inst80 (
                                            .x(m_dec[80]),
                                            .d(16),
                                            .result(decom_out[80])
                                        );
                                        
                                        decompress_module decompress_inst81 (
                                            .x(m_dec[81]),
                                            .d(16),
                                            .result(decom_out[81])
                                        );
                                        
                                        decompress_module decompress_inst82 (
                                            .x(m_dec[82]),
                                            .d(16),
                                            .result(decom_out[82])
                                        );
                                        
                                        decompress_module decompress_inst83 (
                                            .x(m_dec[83]),
                                            .d(16),
                                            .result(decom_out[83])
                                        );
                                        
                                        decompress_module decompress_inst84 (
                                            .x(m_dec[84]),
                                            .d(16),
                                            .result(decom_out[84])
                                        );
                                        
                                        decompress_module decompress_inst85 (
                                            .x(m_dec[85]),
                                            .d(16),
                                            .result(decom_out[85])
                                        );
                                        
                                        decompress_module decompress_inst86 (
                                            .x(m_dec[86]),
                                            .d(16),
                                            .result(decom_out[86])
                                        );
                                        
                                        decompress_module decompress_inst87 (
                                            .x(m_dec[87]),
                                            .d(16),
                                            .result(decom_out[87])
                                        );
                                        
                                        decompress_module decompress_inst88 (
                                            .x(m_dec[88]),
                                            .d(16),
                                            .result(decom_out[88])
                                        );
                                        
                                        decompress_module decompress_inst89 (
                                            .x(m_dec[89]),
                                            .d(16),
                                            .result(decom_out[89])
                                        );
                                        
                                        decompress_module decompress_inst90 (
                                            .x(m_dec[90]),
                                            .d(16),
                                            .result(decom_out[90])
                                        );
                                        
                                        decompress_module decompress_inst91 (
                                            .x(m_dec[91]),
                                            .d(16),
                                            .result(decom_out[91])
                                        );
                                        
                                        decompress_module decompress_inst92 (
                                            .x(m_dec[92]),
                                            .d(16),
                                            .result(decom_out[92])
                                        );
                                        
                                        decompress_module decompress_inst93 (
                                            .x(m_dec[93]),
                                            .d(16),
                                            .result(decom_out[93])
                                        );
                                        
                                        decompress_module decompress_inst94 (
                                            .x(m_dec[94]),
                                            .d(16),
                                            .result(decom_out[94])
                                        );
                                        
                                        decompress_module decompress_inst95 (
                                            .x(m_dec[95]),
                                            .d(16),
                                            .result(decom_out[95])
                                        );
                                        
                                        decompress_module decompress_inst96 (
                                            .x(m_dec[96]),
                                            .d(16),
                                            .result(decom_out[96])
                                        );
                                        
                                        decompress_module decompress_inst97 (
                                            .x(m_dec[97]),
                                            .d(16),
                                            .result(decom_out[97])
                                        );
                                        
                                        decompress_module decompress_inst98 (
                                            .x(m_dec[98]),
                                            .d(16),
                                            .result(decom_out[98])
                                        );
                                        
                                        decompress_module decompress_inst99 (
                                            .x(m_dec[99]),
                                            .d(16),
                                            .result(decom_out[99])
                                        );
                                        
                                        decompress_module decompress_inst100 (
                                            .x(m_dec[100]),
                                            .d(16),
                                            .result(decom_out[100])
                                        );
                                        
                                        decompress_module decompress_inst101 (
                                            .x(m_dec[101]),
                                            .d(16),
                                            .result(decom_out[101])
                                        );
                                        
                                        decompress_module decompress_inst102 (
                                            .x(m_dec[102]),
                                            .d(16),
                                            .result(decom_out[102])
                                        );
                                        
                                        decompress_module decompress_inst103 (
                                            .x(m_dec[103]),
                                            .d(16),
                                            .result(decom_out[103])
                                        );
                                        
                                        decompress_module decompress_inst104 (
                                            .x(m_dec[104]),
                                            .d(16),
                                            .result(decom_out[104])
                                        );
                                        
                                        decompress_module decompress_inst105 (
                                            .x(m_dec[105]),
                                            .d(16),
                                            .result(decom_out[105])
                                        );
                                        
                                        decompress_module decompress_inst106 (
                                            .x(m_dec[106]),
                                            .d(16),
                                            .result(decom_out[106])
                                        );
                                        
                                        decompress_module decompress_inst107 (
                                            .x(m_dec[107]),
                                            .d(16),
                                            .result(decom_out[107])
                                        );
                                        
                                        decompress_module decompress_inst108 (
                                            .x(m_dec[108]),
                                            .d(16),
                                            .result(decom_out[108])
                                        );
                                        
                                        decompress_module decompress_inst109 (
                                            .x(m_dec[109]),
                                            .d(16),
                                            .result(decom_out[109])
                                        );
                                        
                                        decompress_module decompress_inst110 (
                                            .x(m_dec[110]),
                                            .d(16),
                                            .result(decom_out[110])
                                        );
                                        
                                        decompress_module decompress_inst111 (
                                            .x(m_dec[111]),
                                            .d(16),
                                            .result(decom_out[111])
                                        );
                                        
                                        decompress_module decompress_inst112 (
                                            .x(m_dec[112]),
                                            .d(16),
                                            .result(decom_out[112])
                                        );
                                        
                                        decompress_module decompress_inst113 (
                                            .x(m_dec[113]),
                                            .d(16),
                                            .result(decom_out[113])
                                        );
                                        
                                        decompress_module decompress_inst114 (
                                            .x(m_dec[114]),
                                            .d(16),
                                            .result(decom_out[114])
                                        );
                                        
                                        decompress_module decompress_inst115 (
                                            .x(m_dec[115]),
                                            .d(16),
                                            .result(decom_out[115])
                                        );
                                        
                                        decompress_module decompress_inst116 (
                                            .x(m_dec[116]),
                                            .d(16),
                                            .result(decom_out[116])
                                        );
                                        
                                        decompress_module decompress_inst117 (
                                            .x(m_dec[117]),
                                            .d(16),
                                            .result(decom_out[117])
                                        );
                                        
                                        decompress_module decompress_inst118 (
                                            .x(m_dec[118]),
                                            .d(16),
                                            .result(decom_out[118])
                                        );
                                        
                                        decompress_module decompress_inst119 (
                                            .x(m_dec[119]),
                                            .d(16),
                                            .result(decom_out[119])
                                        );
                                        
                                        decompress_module decompress_inst120 (
                                            .x(m_dec[120]),
                                            .d(16),
                                            .result(decom_out[120])
                                        );
                                        
                                        decompress_module decompress_inst121 (
                                            .x(m_dec[121]),
                                            .d(16),
                                            .result(decom_out[121])
                                        );
                                        
                                        decompress_module decompress_inst122 (
                                            .x(m_dec[122]),
                                            .d(16),
                                            .result(decom_out[122])
                                        );
                                        
                                        decompress_module decompress_inst123 (
                                            .x(m_dec[123]),
                                            .d(16),
                                            .result(decom_out[123])
                                        );
                                        
                                        decompress_module decompress_inst124 (
                                            .x(m_dec[124]),
                                            .d(16),
                                            .result(decom_out[124])
                                        );
                                        
                                        decompress_module decompress_inst125 (
                                            .x(m_dec[125]),
                                            .d(16),
                                            .result(decom_out[125])
                                        );
                                        
                                        decompress_module decompress_inst126 (
                                            .x(m_dec[126]),
                                            .d(16),
                                            .result(decom_out[126])
                                        );
                                        
                                        decompress_module decompress_inst127 (
                                            .x(m_dec[127]),
                                            .d(16),
                                            .result(decom_out[127])
                                        );
                                        
                                        decompress_module decompress_inst128 (
                                            .x(m_dec[128]),
                                            .d(16),
                                            .result(decom_out[128])
                                        );
                                        
                                        decompress_module decompress_inst129 (
                                            .x(m_dec[129]),
                                            .d(16),
                                            .result(decom_out[129])
                                        );
                                        
                                        decompress_module decompress_inst130 (
                                            .x(m_dec[130]),
                                            .d(16),
                                            .result(decom_out[130])
                                        );
                                        
                                        decompress_module decompress_inst131 (
                                            .x(m_dec[131]),
                                            .d(16),
                                            .result(decom_out[131])
                                        );
                                        
                                        decompress_module decompress_inst132 (
                                            .x(m_dec[132]),
                                            .d(16),
                                            .result(decom_out[132])
                                        );
                                        
                                        decompress_module decompress_inst133 (
                                            .x(m_dec[133]),
                                            .d(16),
                                            .result(decom_out[133])
                                        );
                                        
                                        decompress_module decompress_inst134 (
                                            .x(m_dec[134]),
                                            .d(16),
                                            .result(decom_out[134])
                                        );
                                        
                                        decompress_module decompress_inst135 (
                                            .x(m_dec[135]),
                                            .d(16),
                                            .result(decom_out[135])
                                        );
                                        
                                        decompress_module decompress_inst136 (
                                            .x(m_dec[136]),
                                            .d(16),
                                            .result(decom_out[136])
                                        );
                                        
                                        decompress_module decompress_inst137 (
                                            .x(m_dec[137]),
                                            .d(16),
                                            .result(decom_out[137])
                                        );
                                        
                                        decompress_module decompress_inst138 (
                                            .x(m_dec[138]),
                                            .d(16),
                                            .result(decom_out[138])
                                        );
                                        
                                        decompress_module decompress_inst139 (
                                            .x(m_dec[139]),
                                            .d(16),
                                            .result(decom_out[139])
                                        );
                                        
                                        decompress_module decompress_inst140 (
                                            .x(m_dec[140]),
                                            .d(16),
                                            .result(decom_out[140])
                                        );
                                        
                                        decompress_module decompress_inst141 (
                                            .x(m_dec[141]),
                                            .d(16),
                                            .result(decom_out[141])
                                        );
                                        
                                        decompress_module decompress_inst142 (
                                            .x(m_dec[142]),
                                            .d(16),
                                            .result(decom_out[142])
                                        );
                                        
                                        decompress_module decompress_inst143 (
                                            .x(m_dec[143]),
                                            .d(16),
                                            .result(decom_out[143])
                                        );
                                        
                                        decompress_module decompress_inst144 (
                                            .x(m_dec[144]),
                                            .d(16),
                                            .result(decom_out[144])
                                        );
                                        
                                        decompress_module decompress_inst145 (
                                            .x(m_dec[145]),
                                            .d(16),
                                            .result(decom_out[145])
                                        );
                                        
                                        decompress_module decompress_inst146 (
                                            .x(m_dec[146]),
                                            .d(16),
                                            .result(decom_out[146])
                                        );
                                        
                                        decompress_module decompress_inst147 (
                                            .x(m_dec[147]),
                                            .d(16),
                                            .result(decom_out[147])
                                        );
                                        
                                        decompress_module decompress_inst148 (
                                            .x(m_dec[148]),
                                            .d(16),
                                            .result(decom_out[148])
                                        );
                                        
                                        decompress_module decompress_inst149 (
                                            .x(m_dec[149]),
                                            .d(16),
                                            .result(decom_out[149])
                                        );
                                        
                                        decompress_module decompress_inst150 (
                                            .x(m_dec[150]),
                                            .d(16),
                                            .result(decom_out[150])
                                        );
                                        
                                        decompress_module decompress_inst151 (
                                            .x(m_dec[151]),
                                            .d(16),
                                            .result(decom_out[151])
                                        );
                                        
                                        decompress_module decompress_inst152 (
                                            .x(m_dec[152]),
                                            .d(16),
                                            .result(decom_out[152])
                                        );
                                        
                                        decompress_module decompress_inst153 (
                                            .x(m_dec[153]),
                                            .d(16),
                                            .result(decom_out[153])
                                        );
                                        
                                        decompress_module decompress_inst154 (
                                            .x(m_dec[154]),
                                            .d(16),
                                            .result(decom_out[154])
                                        );
                                        
                                        decompress_module decompress_inst155 (
                                            .x(m_dec[155]),
                                            .d(16),
                                            .result(decom_out[155])
                                        );
                                        
                                        decompress_module decompress_inst156 (
                                            .x(m_dec[156]),
                                            .d(16),
                                            .result(decom_out[156])
                                        );
                                        
                                        decompress_module decompress_inst157 (
                                            .x(m_dec[157]),
                                            .d(16),
                                            .result(decom_out[157])
                                        );
                                        
                                        decompress_module decompress_inst158 (
                                            .x(m_dec[158]),
                                            .d(16),
                                            .result(decom_out[158])
                                        );
                                        
                                        decompress_module decompress_inst159 (
                                            .x(m_dec[159]),
                                            .d(16),
                                            .result(decom_out[159])
                                        );
                                        
                                        decompress_module decompress_inst160 (
                                            .x(m_dec[160]),
                                            .d(16),
                                            .result(decom_out[160])
                                        );
                                        
                                        decompress_module decompress_inst161 (
                                            .x(m_dec[161]),
                                            .d(16),
                                            .result(decom_out[161])
                                        );
                                        
                                        decompress_module decompress_inst162 (
                                            .x(m_dec[162]),
                                            .d(16),
                                            .result(decom_out[162])
                                        );
                                        
                                        decompress_module decompress_inst163 (
                                            .x(m_dec[163]),
                                            .d(16),
                                            .result(decom_out[163])
                                        );
                                        
                                        decompress_module decompress_inst164 (
                                            .x(m_dec[164]),
                                            .d(16),
                                            .result(decom_out[164])
                                        );
                                        
                                        decompress_module decompress_inst165 (
                                            .x(m_dec[165]),
                                            .d(16),
                                            .result(decom_out[165])
                                        );
                                        
                                        decompress_module decompress_inst166 (
                                            .x(m_dec[166]),
                                            .d(16),
                                            .result(decom_out[166])
                                        );
                                        
                                        decompress_module decompress_inst167 (
                                            .x(m_dec[167]),
                                            .d(16),
                                            .result(decom_out[167])
                                        );
                                        
                                        decompress_module decompress_inst168 (
                                            .x(m_dec[168]),
                                            .d(16),
                                            .result(decom_out[168])
                                        );
                                        
                                        decompress_module decompress_inst169 (
                                            .x(m_dec[169]),
                                            .d(16),
                                            .result(decom_out[169])
                                        );
                                        
                                        decompress_module decompress_inst170 (
                                            .x(m_dec[170]),
                                            .d(16),
                                            .result(decom_out[170])
                                        );
                                        
                                        decompress_module decompress_inst171 (
                                            .x(m_dec[171]),
                                            .d(16),
                                            .result(decom_out[171])
                                        );
                                        
                                        decompress_module decompress_inst172 (
                                            .x(m_dec[172]),
                                            .d(16),
                                            .result(decom_out[172])
                                        );
                                        
                                        decompress_module decompress_inst173 (
                                            .x(m_dec[173]),
                                            .d(16),
                                            .result(decom_out[173])
                                        );
                                        
                                        decompress_module decompress_inst174 (
                                            .x(m_dec[174]),
                                            .d(16),
                                            .result(decom_out[174])
                                        );
                                        
                                        decompress_module decompress_inst175 (
                                            .x(m_dec[175]),
                                            .d(16),
                                            .result(decom_out[175])
                                        );
                                        
                                        decompress_module decompress_inst176 (
                                            .x(m_dec[176]),
                                            .d(16),
                                            .result(decom_out[176])
                                        );
                                        
                                        decompress_module decompress_inst177 (
                                            .x(m_dec[177]),
                                            .d(16),
                                            .result(decom_out[177])
                                        );
                                        
                                        decompress_module decompress_inst178 (
                                            .x(m_dec[178]),
                                            .d(16),
                                            .result(decom_out[178])
                                        );
                                        
                                        decompress_module decompress_inst179 (
                                            .x(m_dec[179]),
                                            .d(16),
                                            .result(decom_out[179])
                                        );
                                        
                                        decompress_module decompress_inst180 (
                                            .x(m_dec[180]),
                                            .d(16),
                                            .result(decom_out[180])
                                        );
                                        
                                        decompress_module decompress_inst181 (
                                            .x(m_dec[181]),
                                            .d(16),
                                            .result(decom_out[181])
                                        );
                                        
                                        decompress_module decompress_inst182 (
                                            .x(m_dec[182]),
                                            .d(16),
                                            .result(decom_out[182])
                                        );
                                        
                                        decompress_module decompress_inst183 (
                                            .x(m_dec[183]),
                                            .d(16),
                                            .result(decom_out[183])
                                        );
                                        
                                        decompress_module decompress_inst184 (
                                            .x(m_dec[184]),
                                            .d(16),
                                            .result(decom_out[184])
                                        );
                                        
                                        decompress_module decompress_inst185 (
                                            .x(m_dec[185]),
                                            .d(16),
                                            .result(decom_out[185])
                                        );
                                        
                                        decompress_module decompress_inst186 (
                                            .x(m_dec[186]),
                                            .d(16),
                                            .result(decom_out[186])
                                        );
                                        
                                        decompress_module decompress_inst187 (
                                            .x(m_dec[187]),
                                            .d(16),
                                            .result(decom_out[187])
                                        );
                                        
                                        decompress_module decompress_inst188 (
                                            .x(m_dec[188]),
                                            .d(16),
                                            .result(decom_out[188])
                                        );
                                        
                                        decompress_module decompress_inst189 (
                                            .x(m_dec[189]),
                                            .d(16),
                                            .result(decom_out[189])
                                        );
                                        
                                        decompress_module decompress_inst190 (
                                            .x(m_dec[190]),
                                            .d(16),
                                            .result(decom_out[190])
                                        );
                                        
                                        decompress_module decompress_inst191 (
                                            .x(m_dec[191]),
                                            .d(16),
                                            .result(decom_out[191])
                                        );
                                        
                                        decompress_module decompress_inst192 (
                                            .x(m_dec[192]),
                                            .d(16),
                                            .result(decom_out[192])
                                        );
                                        
                                        decompress_module decompress_inst193 (
                                            .x(m_dec[193]),
                                            .d(16),
                                            .result(decom_out[193])
                                        );
                                        
                                        decompress_module decompress_inst194 (
                                            .x(m_dec[194]),
                                            .d(16),
                                            .result(decom_out[194])
                                        );
                                        
                                        decompress_module decompress_inst195 (
                                            .x(m_dec[195]),
                                            .d(16),
                                            .result(decom_out[195])
                                        );
                                        
                                        decompress_module decompress_inst196 (
                                            .x(m_dec[196]),
                                            .d(16),
                                            .result(decom_out[196])
                                        );
                                        
                                        decompress_module decompress_inst197 (
                                            .x(m_dec[197]),
                                            .d(16),
                                            .result(decom_out[197])
                                        );
                                        
                                        decompress_module decompress_inst198 (
                                            .x(m_dec[198]),
                                            .d(16),
                                            .result(decom_out[198])
                                        );
                                        
                                        decompress_module decompress_inst199 (
                                            .x(m_dec[199]),
                                            .d(16),
                                            .result(decom_out[199])
                                        );
                                        
                                        decompress_module decompress_inst200 (
                                            .x(m_dec[200]),
                                            .d(16),
                                            .result(decom_out[200])
                                        );
                                        
                                        decompress_module decompress_inst201 (
                                            .x(m_dec[201]),
                                            .d(16),
                                            .result(decom_out[201])
                                        );
                                        
                                        decompress_module decompress_inst202 (
                                            .x(m_dec[202]),
                                            .d(16),
                                            .result(decom_out[202])
                                        );
                                        
                                        decompress_module decompress_inst203 (
                                            .x(m_dec[203]),
                                            .d(16),
                                            .result(decom_out[203])
                                        );
                                        
                                        decompress_module decompress_inst204 (
                                            .x(m_dec[204]),
                                            .d(16),
                                            .result(decom_out[204])
                                        );
                                        
                                        decompress_module decompress_inst205 (
                                            .x(m_dec[205]),
                                            .d(16),
                                            .result(decom_out[205])
                                        );
                                        
                                        decompress_module decompress_inst206 (
                                            .x(m_dec[206]),
                                            .d(16),
                                            .result(decom_out[206])
                                        );
                                        
                                        decompress_module decompress_inst207 (
                                            .x(m_dec[207]),
                                            .d(16),
                                            .result(decom_out[207])
                                        );
                                        
                                        decompress_module decompress_inst208 (
                                            .x(m_dec[208]),
                                            .d(16),
                                            .result(decom_out[208])
                                        );
                                        
                                        decompress_module decompress_inst209 (
                                            .x(m_dec[209]),
                                            .d(16),
                                            .result(decom_out[209])
                                        );
                                        
                                        decompress_module decompress_inst210 (
                                            .x(m_dec[210]),
                                            .d(16),
                                            .result(decom_out[210])
                                        );
                                        
                                        decompress_module decompress_inst211 (
                                            .x(m_dec[211]),
                                            .d(16),
                                            .result(decom_out[211])
                                        );
                                        
                                        decompress_module decompress_inst212 (
                                            .x(m_dec[212]),
                                            .d(16),
                                            .result(decom_out[212])
                                        );
                                        
                                        decompress_module decompress_inst213 (
                                            .x(m_dec[213]),
                                            .d(16),
                                            .result(decom_out[213])
                                        );
                                        
                                        decompress_module decompress_inst214 (
                                            .x(m_dec[214]),
                                            .d(16),
                                            .result(decom_out[214])
                                        );
                                        
                                        decompress_module decompress_inst215 (
                                            .x(m_dec[215]),
                                            .d(16),
                                            .result(decom_out[215])
                                        );
                                        
                                        decompress_module decompress_inst216 (
                                            .x(m_dec[216]),
                                            .d(16),
                                            .result(decom_out[216])
                                        );
                                        
                                        decompress_module decompress_inst217 (
                                            .x(m_dec[217]),
                                            .d(16),
                                            .result(decom_out[217])
                                        );
                                        
                                        decompress_module decompress_inst218 (
                                            .x(m_dec[218]),
                                            .d(16),
                                            .result(decom_out[218])
                                        );
                                        
                                        decompress_module decompress_inst219 (
                                            .x(m_dec[219]),
                                            .d(16),
                                            .result(decom_out[219])
                                        );
                                        
                                        decompress_module decompress_inst220 (
                                            .x(m_dec[220]),
                                            .d(16),
                                            .result(decom_out[220])
                                        );
                                        
                                        decompress_module decompress_inst221 (
                                            .x(m_dec[221]),
                                            .d(16),
                                            .result(decom_out[221])
                                        );
                                        
                                        decompress_module decompress_inst222 (
                                            .x(m_dec[222]),
                                            .d(16),
                                            .result(decom_out[222])
                                        );
                                        
                                        decompress_module decompress_inst223 (
                                            .x(m_dec[223]),
                                            .d(16),
                                            .result(decom_out[223])
                                        );
                                        
                                        decompress_module decompress_inst224 (
                                            .x(m_dec[224]),
                                            .d(16),
                                            .result(decom_out[224])
                                        );
                                        
                                        decompress_module decompress_inst225 (
                                            .x(m_dec[225]),
                                            .d(16),
                                            .result(decom_out[225])
                                        );
                                        
                                        decompress_module decompress_inst226 (
                                            .x(m_dec[226]),
                                            .d(16),
                                            .result(decom_out[226])
                                        );
                                        
                                        decompress_module decompress_inst227 (
                                            .x(m_dec[227]),
                                            .d(16),
                                            .result(decom_out[227])
                                        );
                                        
                                        decompress_module decompress_inst228 (
                                            .x(m_dec[228]),
                                            .d(16),
                                            .result(decom_out[228])
                                        );
                                        
                                        decompress_module decompress_inst229 (
                                            .x(m_dec[229]),
                                            .d(16),
                                            .result(decom_out[229])
                                        );
                                        
                                        decompress_module decompress_inst230 (
                                            .x(m_dec[230]),
                                            .d(16),
                                            .result(decom_out[230])
                                        );
                                        
                                        decompress_module decompress_inst231 (
                                            .x(m_dec[231]),
                                            .d(16),
                                            .result(decom_out[231])
                                        );
                                        
                                        decompress_module decompress_inst232 (
                                            .x(m_dec[232]),
                                            .d(16),
                                            .result(decom_out[232])
                                        );
                                        
                                        decompress_module decompress_inst233 (
                                            .x(m_dec[233]),
                                            .d(16),
                                            .result(decom_out[233])
                                        );
                                        
                                        decompress_module decompress_inst234 (
                                            .x(m_dec[234]),
                                            .d(16),
                                            .result(decom_out[234])
                                        );
                                        
                                        decompress_module decompress_inst235 (
                                            .x(m_dec[235]),
                                            .d(16),
                                            .result(decom_out[235])
                                        );
                                        
                                        decompress_module decompress_inst236 (
                                            .x(m_dec[236]),
                                            .d(16),
                                            .result(decom_out[236])
                                        );
                                        
                                        decompress_module decompress_inst237 (
                                            .x(m_dec[237]),
                                            .d(16),
                                            .result(decom_out[237])
                                        );
                                        
                                        decompress_module decompress_inst238 (
                                            .x(m_dec[238]),
                                            .d(16),
                                            .result(decom_out[238])
                                        );
                                        
                                        decompress_module decompress_inst239 (
                                            .x(m_dec[239]),
                                            .d(16),
                                            .result(decom_out[239])
                                        );
                                        
                                        decompress_module decompress_inst240 (
                                            .x(m_dec[240]),
                                            .d(16),
                                            .result(decom_out[240])
                                        );
                                        
                                        decompress_module decompress_inst241 (
                                            .x(m_dec[241]),
                                            .d(16),
                                            .result(decom_out[241])
                                        );
                                        
                                        decompress_module decompress_inst242 (
                                            .x(m_dec[242]),
                                            .d(16),
                                            .result(decom_out[242])
                                        );
                                        
                                        decompress_module decompress_inst243 (
                                            .x(m_dec[243]),
                                            .d(16),
                                            .result(decom_out[243])
                                        );
                                        
                                        decompress_module decompress_inst244 (
                                            .x(m_dec[244]),
                                            .d(16),
                                            .result(decom_out[244])
                                        );
                                        
                                        decompress_module decompress_inst245 (
                                            .x(m_dec[245]),
                                            .d(16),
                                            .result(decom_out[245])
                                        );
                                        
                                        decompress_module decompress_inst246 (
                                            .x(m_dec[246]),
                                            .d(16),
                                            .result(decom_out[246])
                                        );
                                        
                                        decompress_module decompress_inst247 (
                                            .x(m_dec[247]),
                                            .d(16),
                                            .result(decom_out[247])
                                        );
                                        
                                        decompress_module decompress_inst248 (
                                            .x(m_dec[248]),
                                            .d(16),
                                            .result(decom_out[248])
                                        );
                                        
                                        decompress_module decompress_inst249 (
                                            .x(m_dec[249]),
                                            .d(16),
                                            .result(decom_out[249])
                                        );
                                        
                                        decompress_module decompress_inst250 (
                                            .x(m_dec[250]),
                                            .d(16),
                                            .result(decom_out[250])
                                        );
                                        
                                        decompress_module decompress_inst251 (
                                            .x(m_dec[251]),
                                            .d(16),
                                            .result(decom_out[251])
                                        );
                                        
                                        decompress_module decompress_inst252 (
                                            .x(m_dec[252]),
                                            .d(16),
                                            .result(decom_out[252])
                                        );
                                        
                                        decompress_module decompress_inst253 (
                                            .x(m_dec[253]),
                                            .d(16),
                                            .result(decom_out[253])
                                        );
                                        
                                        decompress_module decompress_inst254 (
                                            .x(m_dec[254]),
                                            .d(16),
                                            .result(decom_out[254])
                                        );
                                        
                                        decompress_module decompress_inst255 (
                                            .x(m_dec[255]),
                                            .d(16),
                                            .result(decom_out[255])
                                        );
                                        compress_module compress_0 (
                                            .x(u[0][0]),
                                            .d(10),
                                            .result(com_out[0][0])
                                        );
                                        
                                        compress_module compress_1 (
                                            .x(u[0][1]),
                                            .d(10),
                                            .result(com_out[0][1])
                                        );
                                        
                                        compress_module compress_2 (
                                            .x(u[0][2]),
                                            .d(10),
                                            .result(com_out[0][2])
                                        );
                                        
                                        compress_module compress_3 (
                                            .x(u[0][3]),
                                            .d(10),
                                            .result(com_out[0][3])
                                        );
                                        
                                        compress_module compress_4 (
                                            .x(u[0][4]),
                                            .d(10),
                                            .result(com_out[0][4])
                                        );
                                        
                                        compress_module compress_5 (
                                            .x(u[0][5]),
                                            .d(10),
                                            .result(com_out[0][5])
                                        );
                                        
                                        compress_module compress_6 (
                                            .x(u[0][6]),
                                            .d(10),
                                            .result(com_out[0][6])
                                        );
                                        
                                        compress_module compress_7 (
                                            .x(u[0][7]),
                                            .d(10),
                                            .result(com_out[0][7])
                                        );
                                        
                                        compress_module compress_8 (
                                            .x(u[0][8]),
                                            .d(10),
                                            .result(com_out[0][8])
                                        );
                                        
                                        compress_module compress_9 (
                                            .x(u[0][9]),
                                            .d(10),
                                            .result(com_out[0][9])
                                        );
                                        
                                        compress_module compress_10 (
                                            .x(u[0][10]),
                                            .d(10),
                                            .result(com_out[0][10])
                                        );
                                        
                                        compress_module compress_11 (
                                            .x(u[0][11]),
                                            .d(10),
                                            .result(com_out[0][11])
                                        );
                                        
                                        compress_module compress_12 (
                                            .x(u[0][12]),
                                            .d(10),
                                            .result(com_out[0][12])
                                        );
                                        
                                        compress_module compress_13 (
                                            .x(u[0][13]),
                                            .d(10),
                                            .result(com_out[0][13])
                                        );
                                        
                                        compress_module compress_14 (
                                            .x(u[0][14]),
                                            .d(10),
                                            .result(com_out[0][14])
                                        );
                                        
                                        compress_module compress_15 (
                                            .x(u[0][15]),
                                            .d(10),
                                            .result(com_out[0][15])
                                        );
                                        
                                        compress_module compress_16 (
                                            .x(u[0][16]),
                                            .d(10),
                                            .result(com_out[0][16])
                                        );
                                        
                                        compress_module compress_17 (
                                            .x(u[0][17]),
                                            .d(10),
                                            .result(com_out[0][17])
                                        );
                                        
                                        compress_module compress_18 (
                                            .x(u[0][18]),
                                            .d(10),
                                            .result(com_out[0][18])
                                        );
                                        
                                        compress_module compress_19 (
                                            .x(u[0][19]),
                                            .d(10),
                                            .result(com_out[0][19])
                                        );
                                        
                                        compress_module compress_20 (
                                            .x(u[0][20]),
                                            .d(10),
                                            .result(com_out[0][20])
                                        );
                                        
                                        compress_module compress_21 (
                                            .x(u[0][21]),
                                            .d(10),
                                            .result(com_out[0][21])
                                        );
                                        
                                        compress_module compress_22 (
                                            .x(u[0][22]),
                                            .d(10),
                                            .result(com_out[0][22])
                                        );
                                        
                                        compress_module compress_23 (
                                            .x(u[0][23]),
                                            .d(10),
                                            .result(com_out[0][23])
                                        );
                                        
                                        compress_module compress_24 (
                                            .x(u[0][24]),
                                            .d(10),
                                            .result(com_out[0][24])
                                        );
                                        
                                        compress_module compress_25 (
                                            .x(u[0][25]),
                                            .d(10),
                                            .result(com_out[0][25])
                                        );
                                        
                                        compress_module compress_26 (
                                            .x(u[0][26]),
                                            .d(10),
                                            .result(com_out[0][26])
                                        );
                                        
                                        compress_module compress_27 (
                                            .x(u[0][27]),
                                            .d(10),
                                            .result(com_out[0][27])
                                        );
                                        
                                        compress_module compress_28 (
                                            .x(u[0][28]),
                                            .d(10),
                                            .result(com_out[0][28])
                                        );
                                        
                                        compress_module compress_29 (
                                            .x(u[0][29]),
                                            .d(10),
                                            .result(com_out[0][29])
                                        );
                                        
                                        compress_module compress_30 (
                                            .x(u[0][30]),
                                            .d(10),
                                            .result(com_out[0][30])
                                        );
                                        
                                        compress_module compress_31 (
                                            .x(u[0][31]),
                                            .d(10),
                                            .result(com_out[0][31])
                                        );
                                        
                                        compress_module compress_32 (
                                            .x(u[0][32]),
                                            .d(10),
                                            .result(com_out[0][32])
                                        );
                                        
                                        compress_module compress_33 (
                                            .x(u[0][33]),
                                            .d(10),
                                            .result(com_out[0][33])
                                        );
                                        
                                        compress_module compress_34 (
                                            .x(u[0][34]),
                                            .d(10),
                                            .result(com_out[0][34])
                                        );
                                        
                                        compress_module compress_35 (
                                            .x(u[0][35]),
                                            .d(10),
                                            .result(com_out[0][35])
                                        );
                                        
                                        compress_module compress_36 (
                                            .x(u[0][36]),
                                            .d(10),
                                            .result(com_out[0][36])
                                        );
                                        
                                        compress_module compress_37 (
                                            .x(u[0][37]),
                                            .d(10),
                                            .result(com_out[0][37])
                                        );
                                        
                                        compress_module compress_38 (
                                            .x(u[0][38]),
                                            .d(10),
                                            .result(com_out[0][38])
                                        );
                                        
                                        compress_module compress_39 (
                                            .x(u[0][39]),
                                            .d(10),
                                            .result(com_out[0][39])
                                        );
                                        
                                        compress_module compress_40 (
                                            .x(u[0][40]),
                                            .d(10),
                                            .result(com_out[0][40])
                                        );
                                        
                                        compress_module compress_41 (
                                            .x(u[0][41]),
                                            .d(10),
                                            .result(com_out[0][41])
                                        );
                                        
                                        compress_module compress_42 (
                                            .x(u[0][42]),
                                            .d(10),
                                            .result(com_out[0][42])
                                        );
                                        
                                        compress_module compress_43 (
                                            .x(u[0][43]),
                                            .d(10),
                                            .result(com_out[0][43])
                                        );
                                        
                                        compress_module compress_44 (
                                            .x(u[0][44]),
                                            .d(10),
                                            .result(com_out[0][44])
                                        );
                                        
                                        compress_module compress_45 (
                                            .x(u[0][45]),
                                            .d(10),
                                            .result(com_out[0][45])
                                        );
                                        
                                        compress_module compress_46 (
                                            .x(u[0][46]),
                                            .d(10),
                                            .result(com_out[0][46])
                                        );
                                        
                                        compress_module compress_47 (
                                            .x(u[0][47]),
                                            .d(10),
                                            .result(com_out[0][47])
                                        );
                                        
                                        compress_module compress_48 (
                                            .x(u[0][48]),
                                            .d(10),
                                            .result(com_out[0][48])
                                        );
                                        
                                        compress_module compress_49 (
                                            .x(u[0][49]),
                                            .d(10),
                                            .result(com_out[0][49])
                                        );
                                        
                                        compress_module compress_50 (
                                            .x(u[0][50]),
                                            .d(10),
                                            .result(com_out[0][50])
                                        );
                                        
                                        compress_module compress_51 (
                                            .x(u[0][51]),
                                            .d(10),
                                            .result(com_out[0][51])
                                        );
                                        
                                        compress_module compress_52 (
                                            .x(u[0][52]),
                                            .d(10),
                                            .result(com_out[0][52])
                                        );
                                        
                                        compress_module compress_53 (
                                            .x(u[0][53]),
                                            .d(10),
                                            .result(com_out[0][53])
                                        );
                                        
                                        compress_module compress_54 (
                                            .x(u[0][54]),
                                            .d(10),
                                            .result(com_out[0][54])
                                        );
                                        
                                        compress_module compress_55 (
                                            .x(u[0][55]),
                                            .d(10),
                                            .result(com_out[0][55])
                                        );
                                        
                                        compress_module compress_56 (
                                            .x(u[0][56]),
                                            .d(10),
                                            .result(com_out[0][56])
                                        );
                                        
                                        compress_module compress_57 (
                                            .x(u[0][57]),
                                            .d(10),
                                            .result(com_out[0][57])
                                        );
                                        
                                        compress_module compress_58 (
                                            .x(u[0][58]),
                                            .d(10),
                                            .result(com_out[0][58])
                                        );
                                        
                                        compress_module compress_59 (
                                            .x(u[0][59]),
                                            .d(10),
                                            .result(com_out[0][59])
                                        );
                                        
                                        compress_module compress_60 (
                                            .x(u[0][60]),
                                            .d(10),
                                            .result(com_out[0][60])
                                        );
                                        
                                        compress_module compress_61 (
                                            .x(u[0][61]),
                                            .d(10),
                                            .result(com_out[0][61])
                                        );
                                        
                                        compress_module compress_62 (
                                            .x(u[0][62]),
                                            .d(10),
                                            .result(com_out[0][62])
                                        );
                                        
                                        compress_module compress_63 (
                                            .x(u[0][63]),
                                            .d(10),
                                            .result(com_out[0][63])
                                        );
                                        
                                        compress_module compress_64 (
                                            .x(u[0][64]),
                                            .d(10),
                                            .result(com_out[0][64])
                                        );
                                        
                                        compress_module compress_65 (
                                            .x(u[0][65]),
                                            .d(10),
                                            .result(com_out[0][65])
                                        );
                                        
                                        compress_module compress_66 (
                                            .x(u[0][66]),
                                            .d(10),
                                            .result(com_out[0][66])
                                        );
                                        
                                        compress_module compress_67 (
                                            .x(u[0][67]),
                                            .d(10),
                                            .result(com_out[0][67])
                                        );
                                        
                                        compress_module compress_68 (
                                            .x(u[0][68]),
                                            .d(10),
                                            .result(com_out[0][68])
                                        );
                                        
                                        compress_module compress_69 (
                                            .x(u[0][69]),
                                            .d(10),
                                            .result(com_out[0][69])
                                        );
                                        
                                        compress_module compress_70 (
                                            .x(u[0][70]),
                                            .d(10),
                                            .result(com_out[0][70])
                                        );
                                        
                                        compress_module compress_71 (
                                            .x(u[0][71]),
                                            .d(10),
                                            .result(com_out[0][71])
                                        );
                                        
                                        compress_module compress_72 (
                                            .x(u[0][72]),
                                            .d(10),
                                            .result(com_out[0][72])
                                        );
                                        
                                        compress_module compress_73 (
                                            .x(u[0][73]),
                                            .d(10),
                                            .result(com_out[0][73])
                                        );
                                        
                                        compress_module compress_74 (
                                            .x(u[0][74]),
                                            .d(10),
                                            .result(com_out[0][74])
                                        );
                                        
                                        compress_module compress_75 (
                                            .x(u[0][75]),
                                            .d(10),
                                            .result(com_out[0][75])
                                        );
                                        
                                        compress_module compress_76 (
                                            .x(u[0][76]),
                                            .d(10),
                                            .result(com_out[0][76])
                                        );
                                        
                                        compress_module compress_77 (
                                            .x(u[0][77]),
                                            .d(10),
                                            .result(com_out[0][77])
                                        );
                                        
                                        compress_module compress_78 (
                                            .x(u[0][78]),
                                            .d(10),
                                            .result(com_out[0][78])
                                        );
                                        
                                        compress_module compress_79 (
                                            .x(u[0][79]),
                                            .d(10),
                                            .result(com_out[0][79])
                                        );
                                        
                                        compress_module compress_80 (
                                            .x(u[0][80]),
                                            .d(10),
                                            .result(com_out[0][80])
                                        );
                                        
                                        compress_module compress_81 (
                                            .x(u[0][81]),
                                            .d(10),
                                            .result(com_out[0][81])
                                        );
                                        
                                        compress_module compress_82 (
                                            .x(u[0][82]),
                                            .d(10),
                                            .result(com_out[0][82])
                                        );
                                        
                                        compress_module compress_83 (
                                            .x(u[0][83]),
                                            .d(10),
                                            .result(com_out[0][83])
                                        );
                                        
                                        compress_module compress_84 (
                                            .x(u[0][84]),
                                            .d(10),
                                            .result(com_out[0][84])
                                        );
                                        
                                        compress_module compress_85 (
                                            .x(u[0][85]),
                                            .d(10),
                                            .result(com_out[0][85])
                                        );
                                        
                                        compress_module compress_86 (
                                            .x(u[0][86]),
                                            .d(10),
                                            .result(com_out[0][86])
                                        );
                                        
                                        compress_module compress_87 (
                                            .x(u[0][87]),
                                            .d(10),
                                            .result(com_out[0][87])
                                        );
                                        
                                        compress_module compress_88 (
                                            .x(u[0][88]),
                                            .d(10),
                                            .result(com_out[0][88])
                                        );
                                        
                                        compress_module compress_89 (
                                            .x(u[0][89]),
                                            .d(10),
                                            .result(com_out[0][89])
                                        );
                                        
                                        compress_module compress_90 (
                                            .x(u[0][90]),
                                            .d(10),
                                            .result(com_out[0][90])
                                        );
                                        
                                        compress_module compress_91 (
                                            .x(u[0][91]),
                                            .d(10),
                                            .result(com_out[0][91])
                                        );
                                        
                                        compress_module compress_92 (
                                            .x(u[0][92]),
                                            .d(10),
                                            .result(com_out[0][92])
                                        );
                                        
                                        compress_module compress_93 (
                                            .x(u[0][93]),
                                            .d(10),
                                            .result(com_out[0][93])
                                        );
                                        
                                        compress_module compress_94 (
                                            .x(u[0][94]),
                                            .d(10),
                                            .result(com_out[0][94])
                                        );
                                        
                                        compress_module compress_95 (
                                            .x(u[0][95]),
                                            .d(10),
                                            .result(com_out[0][95])
                                        );
                                        
                                        compress_module compress_96 (
                                            .x(u[0][96]),
                                            .d(10),
                                            .result(com_out[0][96])
                                        );
                                        
                                        compress_module compress_97 (
                                            .x(u[0][97]),
                                            .d(10),
                                            .result(com_out[0][97])
                                        );
                                        
                                        compress_module compress_98 (
                                            .x(u[0][98]),
                                            .d(10),
                                            .result(com_out[0][98])
                                        );
                                        
                                        compress_module compress_99 (
                                            .x(u[0][99]),
                                            .d(10),
                                            .result(com_out[0][99])
                                        );
                                        
                                        compress_module compress_100 (
                                            .x(u[0][100]),
                                            .d(10),
                                            .result(com_out[0][100])
                                        );
                                        
                                        compress_module compress_101 (
                                            .x(u[0][101]),
                                            .d(10),
                                            .result(com_out[0][101])
                                        );
                                        
                                        compress_module compress_102 (
                                            .x(u[0][102]),
                                            .d(10),
                                            .result(com_out[0][102])
                                        );
                                        
                                        compress_module compress_103 (
                                            .x(u[0][103]),
                                            .d(10),
                                            .result(com_out[0][103])
                                        );
                                        
                                        compress_module compress_104 (
                                            .x(u[0][104]),
                                            .d(10),
                                            .result(com_out[0][104])
                                        );
                                        
                                        compress_module compress_105 (
                                            .x(u[0][105]),
                                            .d(10),
                                            .result(com_out[0][105])
                                        );
                                        
                                        compress_module compress_106 (
                                            .x(u[0][106]),
                                            .d(10),
                                            .result(com_out[0][106])
                                        );
                                        
                                        compress_module compress_107 (
                                            .x(u[0][107]),
                                            .d(10),
                                            .result(com_out[0][107])
                                        );
                                        
                                        compress_module compress_108 (
                                            .x(u[0][108]),
                                            .d(10),
                                            .result(com_out[0][108])
                                        );
                                        
                                        compress_module compress_109 (
                                            .x(u[0][109]),
                                            .d(10),
                                            .result(com_out[0][109])
                                        );
                                        
                                        compress_module compress_110 (
                                            .x(u[0][110]),
                                            .d(10),
                                            .result(com_out[0][110])
                                        );
                                        
                                        compress_module compress_111 (
                                            .x(u[0][111]),
                                            .d(10),
                                            .result(com_out[0][111])
                                        );
                                        
                                        compress_module compress_112 (
                                            .x(u[0][112]),
                                            .d(10),
                                            .result(com_out[0][112])
                                        );
                                        
                                        compress_module compress_113 (
                                            .x(u[0][113]),
                                            .d(10),
                                            .result(com_out[0][113])
                                        );
                                        
                                        compress_module compress_114 (
                                            .x(u[0][114]),
                                            .d(10),
                                            .result(com_out[0][114])
                                        );
                                        
                                        compress_module compress_115 (
                                            .x(u[0][115]),
                                            .d(10),
                                            .result(com_out[0][115])
                                        );
                                        
                                        compress_module compress_116 (
                                            .x(u[0][116]),
                                            .d(10),
                                            .result(com_out[0][116])
                                        );
                                        
                                        compress_module compress_117 (
                                            .x(u[0][117]),
                                            .d(10),
                                            .result(com_out[0][117])
                                        );
                                        
                                        compress_module compress_118 (
                                            .x(u[0][118]),
                                            .d(10),
                                            .result(com_out[0][118])
                                        );
                                        
                                        compress_module compress_119 (
                                            .x(u[0][119]),
                                            .d(10),
                                            .result(com_out[0][119])
                                        );
                                        
                                        compress_module compress_120 (
                                            .x(u[0][120]),
                                            .d(10),
                                            .result(com_out[0][120])
                                        );
                                        
                                        compress_module compress_121 (
                                            .x(u[0][121]),
                                            .d(10),
                                            .result(com_out[0][121])
                                        );
                                        
                                        compress_module compress_122 (
                                            .x(u[0][122]),
                                            .d(10),
                                            .result(com_out[0][122])
                                        );
                                        
                                        compress_module compress_123 (
                                            .x(u[0][123]),
                                            .d(10),
                                            .result(com_out[0][123])
                                        );
                                        
                                        compress_module compress_124 (
                                            .x(u[0][124]),
                                            .d(10),
                                            .result(com_out[0][124])
                                        );
                                        
                                        compress_module compress_125 (
                                            .x(u[0][125]),
                                            .d(10),
                                            .result(com_out[0][125])
                                        );
                                        
                                        compress_module compress_126 (
                                            .x(u[0][126]),
                                            .d(10),
                                            .result(com_out[0][126])
                                        );
                                        
                                        compress_module compress_127 (
                                            .x(u[0][127]),
                                            .d(10),
                                            .result(com_out[0][127])
                                        );
                                        
                                        compress_module compress_128 (
                                            .x(u[0][128]),
                                            .d(10),
                                            .result(com_out[0][128])
                                        );
                                        
                                        compress_module compress_129 (
                                            .x(u[0][129]),
                                            .d(10),
                                            .result(com_out[0][129])
                                        );
                                        
                                        compress_module compress_130 (
                                            .x(u[0][130]),
                                            .d(10),
                                            .result(com_out[0][130])
                                        );
                                        
                                        compress_module compress_131 (
                                            .x(u[0][131]),
                                            .d(10),
                                            .result(com_out[0][131])
                                        );
                                        
                                        compress_module compress_132 (
                                            .x(u[0][132]),
                                            .d(10),
                                            .result(com_out[0][132])
                                        );
                                        
                                        compress_module compress_133 (
                                            .x(u[0][133]),
                                            .d(10),
                                            .result(com_out[0][133])
                                        );
                                        
                                        compress_module compress_134 (
                                            .x(u[0][134]),
                                            .d(10),
                                            .result(com_out[0][134])
                                        );
                                        
                                        compress_module compress_135 (
                                            .x(u[0][135]),
                                            .d(10),
                                            .result(com_out[0][135])
                                        );
                                        
                                        compress_module compress_136 (
                                            .x(u[0][136]),
                                            .d(10),
                                            .result(com_out[0][136])
                                        );
                                        
                                        compress_module compress_137 (
                                            .x(u[0][137]),
                                            .d(10),
                                            .result(com_out[0][137])
                                        );
                                        
                                        compress_module compress_138 (
                                            .x(u[0][138]),
                                            .d(10),
                                            .result(com_out[0][138])
                                        );
                                        
                                        compress_module compress_139 (
                                            .x(u[0][139]),
                                            .d(10),
                                            .result(com_out[0][139])
                                        );
                                        
                                        compress_module compress_140 (
                                            .x(u[0][140]),
                                            .d(10),
                                            .result(com_out[0][140])
                                        );
                                        
                                        compress_module compress_141 (
                                            .x(u[0][141]),
                                            .d(10),
                                            .result(com_out[0][141])
                                        );
                                        
                                        compress_module compress_142 (
                                            .x(u[0][142]),
                                            .d(10),
                                            .result(com_out[0][142])
                                        );
                                        
                                        compress_module compress_143 (
                                            .x(u[0][143]),
                                            .d(10),
                                            .result(com_out[0][143])
                                        );
                                        
                                        compress_module compress_144 (
                                            .x(u[0][144]),
                                            .d(10),
                                            .result(com_out[0][144])
                                        );
                                        
                                        compress_module compress_145 (
                                            .x(u[0][145]),
                                            .d(10),
                                            .result(com_out[0][145])
                                        );
                                        
                                        compress_module compress_146 (
                                            .x(u[0][146]),
                                            .d(10),
                                            .result(com_out[0][146])
                                        );
                                        
                                        compress_module compress_147 (
                                            .x(u[0][147]),
                                            .d(10),
                                            .result(com_out[0][147])
                                        );
                                        
                                        compress_module compress_148 (
                                            .x(u[0][148]),
                                            .d(10),
                                            .result(com_out[0][148])
                                        );
                                        
                                        compress_module compress_149 (
                                            .x(u[0][149]),
                                            .d(10),
                                            .result(com_out[0][149])
                                        );
                                        
                                        compress_module compress_150 (
                                            .x(u[0][150]),
                                            .d(10),
                                            .result(com_out[0][150])
                                        );
                                        
                                        compress_module compress_151 (
                                            .x(u[0][151]),
                                            .d(10),
                                            .result(com_out[0][151])
                                        );
                                        
                                        compress_module compress_152 (
                                            .x(u[0][152]),
                                            .d(10),
                                            .result(com_out[0][152])
                                        );
                                        
                                        compress_module compress_153 (
                                            .x(u[0][153]),
                                            .d(10),
                                            .result(com_out[0][153])
                                        );
                                        
                                        compress_module compress_154 (
                                            .x(u[0][154]),
                                            .d(10),
                                            .result(com_out[0][154])
                                        );
                                        
                                        compress_module compress_155 (
                                            .x(u[0][155]),
                                            .d(10),
                                            .result(com_out[0][155])
                                        );
                                        
                                        compress_module compress_156 (
                                            .x(u[0][156]),
                                            .d(10),
                                            .result(com_out[0][156])
                                        );
                                        
                                        compress_module compress_157 (
                                            .x(u[0][157]),
                                            .d(10),
                                            .result(com_out[0][157])
                                        );
                                        
                                        compress_module compress_158 (
                                            .x(u[0][158]),
                                            .d(10),
                                            .result(com_out[0][158])
                                        );
                                        
                                        compress_module compress_159 (
                                            .x(u[0][159]),
                                            .d(10),
                                            .result(com_out[0][159])
                                        );
                                        
                                        compress_module compress_160 (
                                            .x(u[0][160]),
                                            .d(10),
                                            .result(com_out[0][160])
                                        );
                                        
                                        compress_module compress_161 (
                                            .x(u[0][161]),
                                            .d(10),
                                            .result(com_out[0][161])
                                        );
                                        
                                        compress_module compress_162 (
                                            .x(u[0][162]),
                                            .d(10),
                                            .result(com_out[0][162])
                                        );
                                        
                                        compress_module compress_163 (
                                            .x(u[0][163]),
                                            .d(10),
                                            .result(com_out[0][163])
                                        );
                                        
                                        compress_module compress_164 (
                                            .x(u[0][164]),
                                            .d(10),
                                            .result(com_out[0][164])
                                        );
                                        
                                        compress_module compress_165 (
                                            .x(u[0][165]),
                                            .d(10),
                                            .result(com_out[0][165])
                                        );
                                        
                                        compress_module compress_166 (
                                            .x(u[0][166]),
                                            .d(10),
                                            .result(com_out[0][166])
                                        );
                                        
                                        compress_module compress_167 (
                                            .x(u[0][167]),
                                            .d(10),
                                            .result(com_out[0][167])
                                        );
                                        
                                        compress_module compress_168 (
                                            .x(u[0][168]),
                                            .d(10),
                                            .result(com_out[0][168])
                                        );
                                        
                                        compress_module compress_169 (
                                            .x(u[0][169]),
                                            .d(10),
                                            .result(com_out[0][169])
                                        );
                                        
                                        compress_module compress_170 (
                                            .x(u[0][170]),
                                            .d(10),
                                            .result(com_out[0][170])
                                        );
                                        
                                        compress_module compress_171 (
                                            .x(u[0][171]),
                                            .d(10),
                                            .result(com_out[0][171])
                                        );
                                        
                                        compress_module compress_172 (
                                            .x(u[0][172]),
                                            .d(10),
                                            .result(com_out[0][172])
                                        );
                                        
                                        compress_module compress_173 (
                                            .x(u[0][173]),
                                            .d(10),
                                            .result(com_out[0][173])
                                        );
                                        
                                        compress_module compress_174 (
                                            .x(u[0][174]),
                                            .d(10),
                                            .result(com_out[0][174])
                                        );
                                        
                                        compress_module compress_175 (
                                            .x(u[0][175]),
                                            .d(10),
                                            .result(com_out[0][175])
                                        );
                                        
                                        compress_module compress_176 (
                                            .x(u[0][176]),
                                            .d(10),
                                            .result(com_out[0][176])
                                        );
                                        
                                        compress_module compress_177 (
                                            .x(u[0][177]),
                                            .d(10),
                                            .result(com_out[0][177])
                                        );
                                        
                                        compress_module compress_178 (
                                            .x(u[0][178]),
                                            .d(10),
                                            .result(com_out[0][178])
                                        );
                                        
                                        compress_module compress_179 (
                                            .x(u[0][179]),
                                            .d(10),
                                            .result(com_out[0][179])
                                        );
                                        
                                        compress_module compress_180 (
                                            .x(u[0][180]),
                                            .d(10),
                                            .result(com_out[0][180])
                                        );
                                        
                                        compress_module compress_181 (
                                            .x(u[0][181]),
                                            .d(10),
                                            .result(com_out[0][181])
                                        );
                                        
                                        compress_module compress_182 (
                                            .x(u[0][182]),
                                            .d(10),
                                            .result(com_out[0][182])
                                        );
                                        
                                        compress_module compress_183 (
                                            .x(u[0][183]),
                                            .d(10),
                                            .result(com_out[0][183])
                                        );
                                        
                                        compress_module compress_184 (
                                            .x(u[0][184]),
                                            .d(10),
                                            .result(com_out[0][184])
                                        );
                                        
                                        compress_module compress_185 (
                                            .x(u[0][185]),
                                            .d(10),
                                            .result(com_out[0][185])
                                        );
                                        
                                        compress_module compress_186 (
                                            .x(u[0][186]),
                                            .d(10),
                                            .result(com_out[0][186])
                                        );
                                        
                                        compress_module compress_187 (
                                            .x(u[0][187]),
                                            .d(10),
                                            .result(com_out[0][187])
                                        );
                                        
                                        compress_module compress_188 (
                                            .x(u[0][188]),
                                            .d(10),
                                            .result(com_out[0][188])
                                        );
                                        
                                        compress_module compress_189 (
                                            .x(u[0][189]),
                                            .d(10),
                                            .result(com_out[0][189])
                                        );
                                        
                                        compress_module compress_190 (
                                            .x(u[0][190]),
                                            .d(10),
                                            .result(com_out[0][190])
                                        );
                                        
                                        compress_module compress_191 (
                                            .x(u[0][191]),
                                            .d(10),
                                            .result(com_out[0][191])
                                        );
                                        
                                        compress_module compress_192 (
                                            .x(u[0][192]),
                                            .d(10),
                                            .result(com_out[0][192])
                                        );
                                        
                                        compress_module compress_193 (
                                            .x(u[0][193]),
                                            .d(10),
                                            .result(com_out[0][193])
                                        );
                                        
                                        compress_module compress_194 (
                                            .x(u[0][194]),
                                            .d(10),
                                            .result(com_out[0][194])
                                        );
                                        
                                        compress_module compress_195 (
                                            .x(u[0][195]),
                                            .d(10),
                                            .result(com_out[0][195])
                                        );
                                        
                                        compress_module compress_196 (
                                            .x(u[0][196]),
                                            .d(10),
                                            .result(com_out[0][196])
                                        );
                                        
                                        compress_module compress_197 (
                                            .x(u[0][197]),
                                            .d(10),
                                            .result(com_out[0][197])
                                        );
                                        
                                        compress_module compress_198 (
                                            .x(u[0][198]),
                                            .d(10),
                                            .result(com_out[0][198])
                                        );
                                        
                                        compress_module compress_199 (
                                            .x(u[0][199]),
                                            .d(10),
                                            .result(com_out[0][199])
                                        );
                                        
                                        compress_module compress_200 (
                                            .x(u[0][200]),
                                            .d(10),
                                            .result(com_out[0][200])
                                        );
                                        
                                        compress_module compress_201 (
                                            .x(u[0][201]),
                                            .d(10),
                                            .result(com_out[0][201])
                                        );
                                        
                                        compress_module compress_202 (
                                            .x(u[0][202]),
                                            .d(10),
                                            .result(com_out[0][202])
                                        );
                                        
                                        compress_module compress_203 (
                                            .x(u[0][203]),
                                            .d(10),
                                            .result(com_out[0][203])
                                        );
                                        
                                        compress_module compress_204 (
                                            .x(u[0][204]),
                                            .d(10),
                                            .result(com_out[0][204])
                                        );
                                        
                                        compress_module compress_205 (
                                            .x(u[0][205]),
                                            .d(10),
                                            .result(com_out[0][205])
                                        );
                                        
                                        compress_module compress_206 (
                                            .x(u[0][206]),
                                            .d(10),
                                            .result(com_out[0][206])
                                        );
                                        
                                        compress_module compress_207 (
                                            .x(u[0][207]),
                                            .d(10),
                                            .result(com_out[0][207])
                                        );
                                        
                                        compress_module compress_208 (
                                            .x(u[0][208]),
                                            .d(10),
                                            .result(com_out[0][208])
                                        );
                                        
                                        compress_module compress_209 (
                                            .x(u[0][209]),
                                            .d(10),
                                            .result(com_out[0][209])
                                        );
                                        
                                        compress_module compress_210 (
                                            .x(u[0][210]),
                                            .d(10),
                                            .result(com_out[0][210])
                                        );
                                        
                                        compress_module compress_211 (
                                            .x(u[0][211]),
                                            .d(10),
                                            .result(com_out[0][211])
                                        );
                                        
                                        compress_module compress_212 (
                                            .x(u[0][212]),
                                            .d(10),
                                            .result(com_out[0][212])
                                        );
                                        
                                        compress_module compress_213 (
                                            .x(u[0][213]),
                                            .d(10),
                                            .result(com_out[0][213])
                                        );
                                        
                                        compress_module compress_214 (
                                            .x(u[0][214]),
                                            .d(10),
                                            .result(com_out[0][214])
                                        );
                                        
                                        compress_module compress_215 (
                                            .x(u[0][215]),
                                            .d(10),
                                            .result(com_out[0][215])
                                        );
                                        
                                        compress_module compress_216 (
                                            .x(u[0][216]),
                                            .d(10),
                                            .result(com_out[0][216])
                                        );
                                        
                                        compress_module compress_217 (
                                            .x(u[0][217]),
                                            .d(10),
                                            .result(com_out[0][217])
                                        );
                                        
                                        compress_module compress_218 (
                                            .x(u[0][218]),
                                            .d(10),
                                            .result(com_out[0][218])
                                        );
                                        
                                        compress_module compress_219 (
                                            .x(u[0][219]),
                                            .d(10),
                                            .result(com_out[0][219])
                                        );
                                        
                                        compress_module compress_220 (
                                            .x(u[0][220]),
                                            .d(10),
                                            .result(com_out[0][220])
                                        );
                                        
                                        compress_module compress_221 (
                                            .x(u[0][221]),
                                            .d(10),
                                            .result(com_out[0][221])
                                        );
                                        
                                        compress_module compress_222 (
                                            .x(u[0][222]),
                                            .d(10),
                                            .result(com_out[0][222])
                                        );
                                        
                                        compress_module compress_223 (
                                            .x(u[0][223]),
                                            .d(10),
                                            .result(com_out[0][223])
                                        );
                                        
                                        compress_module compress_224 (
                                            .x(u[0][224]),
                                            .d(10),
                                            .result(com_out[0][224])
                                        );
                                        
                                        compress_module compress_225 (
                                            .x(u[0][225]),
                                            .d(10),
                                            .result(com_out[0][225])
                                        );
                                        
                                        compress_module compress_226 (
                                            .x(u[0][226]),
                                            .d(10),
                                            .result(com_out[0][226])
                                        );
                                        
                                        compress_module compress_227 (
                                            .x(u[0][227]),
                                            .d(10),
                                            .result(com_out[0][227])
                                        );
                                        
                                        compress_module compress_228 (
                                            .x(u[0][228]),
                                            .d(10),
                                            .result(com_out[0][228])
                                        );
                                        
                                        compress_module compress_229 (
                                            .x(u[0][229]),
                                            .d(10),
                                            .result(com_out[0][229])
                                        );
                                        
                                        compress_module compress_230 (
                                            .x(u[0][230]),
                                            .d(10),
                                            .result(com_out[0][230])
                                        );
                                        
                                        compress_module compress_231 (
                                            .x(u[0][231]),
                                            .d(10),
                                            .result(com_out[0][231])
                                        );
                                        
                                        compress_module compress_232 (
                                            .x(u[0][232]),
                                            .d(10),
                                            .result(com_out[0][232])
                                        );
                                        
                                        compress_module compress_233 (
                                            .x(u[0][233]),
                                            .d(10),
                                            .result(com_out[0][233])
                                        );
                                        
                                        compress_module compress_234 (
                                            .x(u[0][234]),
                                            .d(10),
                                            .result(com_out[0][234])
                                        );
                                        
                                        compress_module compress_235 (
                                            .x(u[0][235]),
                                            .d(10),
                                            .result(com_out[0][235])
                                        );
                                        
                                        compress_module compress_236 (
                                            .x(u[0][236]),
                                            .d(10),
                                            .result(com_out[0][236])
                                        );
                                        
                                        compress_module compress_237 (
                                            .x(u[0][237]),
                                            .d(10),
                                            .result(com_out[0][237])
                                        );
                                        
                                        compress_module compress_238 (
                                            .x(u[0][238]),
                                            .d(10),
                                            .result(com_out[0][238])
                                        );
                                        
                                        compress_module compress_239 (
                                            .x(u[0][239]),
                                            .d(10),
                                            .result(com_out[0][239])
                                        );
                                        
                                        compress_module compress_240 (
                                            .x(u[0][240]),
                                            .d(10),
                                            .result(com_out[0][240])
                                        );
                                        
                                        compress_module compress_241 (
                                            .x(u[0][241]),
                                            .d(10),
                                            .result(com_out[0][241])
                                        );
                                        
                                        compress_module compress_242 (
                                            .x(u[0][242]),
                                            .d(10),
                                            .result(com_out[0][242])
                                        );
                                        
                                        compress_module compress_243 (
                                            .x(u[0][243]),
                                            .d(10),
                                            .result(com_out[0][243])
                                        );
                                        
                                        compress_module compress_244 (
                                            .x(u[0][244]),
                                            .d(10),
                                            .result(com_out[0][244])
                                        );
                                        
                                        compress_module compress_245 (
                                            .x(u[0][245]),
                                            .d(10),
                                            .result(com_out[0][245])
                                        );
                                        
                                        compress_module compress_246 (
                                            .x(u[0][246]),
                                            .d(10),
                                            .result(com_out[0][246])
                                        );
                                        
                                        compress_module compress_247 (
                                            .x(u[0][247]),
                                            .d(10),
                                            .result(com_out[0][247])
                                        );
                                        
                                        compress_module compress_248 (
                                            .x(u[0][248]),
                                            .d(10),
                                            .result(com_out[0][248])
                                        );
                                        
                                        compress_module compress_249 (
                                            .x(u[0][249]),
                                            .d(10),
                                            .result(com_out[0][249])
                                        );
                                        
                                        compress_module compress_250 (
                                            .x(u[0][250]),
                                            .d(10),
                                            .result(com_out[0][250])
                                        );
                                        
                                        compress_module compress_251 (
                                            .x(u[0][251]),
                                            .d(10),
                                            .result(com_out[0][251])
                                        );
                                        
                                        compress_module compress_252 (
                                            .x(u[0][252]),
                                            .d(10),
                                            .result(com_out[0][252])
                                        );
                                        
                                        compress_module compress_253 (
                                            .x(u[0][253]),
                                            .d(10),
                                            .result(com_out[0][253])
                                        );
                                        
                                        compress_module compress_254 (
                                            .x(u[0][254]),
                                            .d(10),
                                            .result(com_out[0][254])
                                        );
                                        
                                        compress_module compress_255 (
                                            .x(u[0][255]),
                                            .d(10),
                                            .result(com_out[0][255])
                                        );
                                        
                                        compress_module compress_256 (
                                            .x(u[1][0]),
                                            .d(10),
                                            .result(com_out[1][0])
                                        );
                                        
                                        compress_module compress_257 (
                                            .x(u[1][1]),
                                            .d(10),
                                            .result(com_out[1][1])
                                        );
                                        
                                        compress_module compress_258 (
                                            .x(u[1][2]),
                                            .d(10),
                                            .result(com_out[1][2])
                                        );
                                        
                                        compress_module compress_259 (
                                            .x(u[1][3]),
                                            .d(10),
                                            .result(com_out[1][3])
                                        );
                                        
                                        compress_module compress_260 (
                                            .x(u[1][4]),
                                            .d(10),
                                            .result(com_out[1][4])
                                        );
                                        
                                        compress_module compress_261 (
                                            .x(u[1][5]),
                                            .d(10),
                                            .result(com_out[1][5])
                                        );
                                        
                                        compress_module compress_262 (
                                            .x(u[1][6]),
                                            .d(10),
                                            .result(com_out[1][6])
                                        );
                                        
                                        compress_module compress_263 (
                                            .x(u[1][7]),
                                            .d(10),
                                            .result(com_out[1][7])
                                        );
                                        
                                        compress_module compress_264 (
                                            .x(u[1][8]),
                                            .d(10),
                                            .result(com_out[1][8])
                                        );
                                        
                                        compress_module compress_265 (
                                            .x(u[1][9]),
                                            .d(10),
                                            .result(com_out[1][9])
                                        );
                                        
                                        compress_module compress_266 (
                                            .x(u[1][10]),
                                            .d(10),
                                            .result(com_out[1][10])
                                        );
                                        
                                        compress_module compress_267 (
                                            .x(u[1][11]),
                                            .d(10),
                                            .result(com_out[1][11])
                                        );
                                        
                                        compress_module compress_268 (
                                            .x(u[1][12]),
                                            .d(10),
                                            .result(com_out[1][12])
                                        );
                                        
                                        compress_module compress_269 (
                                            .x(u[1][13]),
                                            .d(10),
                                            .result(com_out[1][13])
                                        );
                                        
                                        compress_module compress_270 (
                                            .x(u[1][14]),
                                            .d(10),
                                            .result(com_out[1][14])
                                        );
                                        
                                        compress_module compress_271 (
                                            .x(u[1][15]),
                                            .d(10),
                                            .result(com_out[1][15])
                                        );
                                        
                                        compress_module compress_272 (
                                            .x(u[1][16]),
                                            .d(10),
                                            .result(com_out[1][16])
                                        );
                                        
                                        compress_module compress_273 (
                                            .x(u[1][17]),
                                            .d(10),
                                            .result(com_out[1][17])
                                        );
                                        
                                        compress_module compress_274 (
                                            .x(u[1][18]),
                                            .d(10),
                                            .result(com_out[1][18])
                                        );
                                        
                                        compress_module compress_275 (
                                            .x(u[1][19]),
                                            .d(10),
                                            .result(com_out[1][19])
                                        );
                                        
                                        compress_module compress_276 (
                                            .x(u[1][20]),
                                            .d(10),
                                            .result(com_out[1][20])
                                        );
                                        
                                        compress_module compress_277 (
                                            .x(u[1][21]),
                                            .d(10),
                                            .result(com_out[1][21])
                                        );
                                        
                                        compress_module compress_278 (
                                            .x(u[1][22]),
                                            .d(10),
                                            .result(com_out[1][22])
                                        );
                                        
                                        compress_module compress_279 (
                                            .x(u[1][23]),
                                            .d(10),
                                            .result(com_out[1][23])
                                        );
                                        
                                        compress_module compress_280 (
                                            .x(u[1][24]),
                                            .d(10),
                                            .result(com_out[1][24])
                                        );
                                        
                                        compress_module compress_281 (
                                            .x(u[1][25]),
                                            .d(10),
                                            .result(com_out[1][25])
                                        );
                                        
                                        compress_module compress_282 (
                                            .x(u[1][26]),
                                            .d(10),
                                            .result(com_out[1][26])
                                        );
                                        
                                        compress_module compress_283 (
                                            .x(u[1][27]),
                                            .d(10),
                                            .result(com_out[1][27])
                                        );
                                        
                                        compress_module compress_284 (
                                            .x(u[1][28]),
                                            .d(10),
                                            .result(com_out[1][28])
                                        );
                                        
                                        compress_module compress_285 (
                                            .x(u[1][29]),
                                            .d(10),
                                            .result(com_out[1][29])
                                        );
                                        
                                        compress_module compress_286 (
                                            .x(u[1][30]),
                                            .d(10),
                                            .result(com_out[1][30])
                                        );
                                        
                                        compress_module compress_287 (
                                            .x(u[1][31]),
                                            .d(10),
                                            .result(com_out[1][31])
                                        );
                                        
                                        compress_module compress_288 (
                                            .x(u[1][32]),
                                            .d(10),
                                            .result(com_out[1][32])
                                        );
                                        
                                        compress_module compress_289 (
                                            .x(u[1][33]),
                                            .d(10),
                                            .result(com_out[1][33])
                                        );
                                        
                                        compress_module compress_290 (
                                            .x(u[1][34]),
                                            .d(10),
                                            .result(com_out[1][34])
                                        );
                                        
                                        compress_module compress_291 (
                                            .x(u[1][35]),
                                            .d(10),
                                            .result(com_out[1][35])
                                        );
                                        
                                        compress_module compress_292 (
                                            .x(u[1][36]),
                                            .d(10),
                                            .result(com_out[1][36])
                                        );
                                        
                                        compress_module compress_293 (
                                            .x(u[1][37]),
                                            .d(10),
                                            .result(com_out[1][37])
                                        );
                                        
                                        compress_module compress_294 (
                                            .x(u[1][38]),
                                            .d(10),
                                            .result(com_out[1][38])
                                        );
                                        
                                        compress_module compress_295 (
                                            .x(u[1][39]),
                                            .d(10),
                                            .result(com_out[1][39])
                                        );
                                        
                                        compress_module compress_296 (
                                            .x(u[1][40]),
                                            .d(10),
                                            .result(com_out[1][40])
                                        );
                                        
                                        compress_module compress_297 (
                                            .x(u[1][41]),
                                            .d(10),
                                            .result(com_out[1][41])
                                        );
                                        
                                        compress_module compress_298 (
                                            .x(u[1][42]),
                                            .d(10),
                                            .result(com_out[1][42])
                                        );
                                        
                                        compress_module compress_299 (
                                            .x(u[1][43]),
                                            .d(10),
                                            .result(com_out[1][43])
                                        );
                                        
                                        compress_module compress_300 (
                                            .x(u[1][44]),
                                            .d(10),
                                            .result(com_out[1][44])
                                        );
                                        
                                        compress_module compress_301 (
                                            .x(u[1][45]),
                                            .d(10),
                                            .result(com_out[1][45])
                                        );
                                        
                                        compress_module compress_302 (
                                            .x(u[1][46]),
                                            .d(10),
                                            .result(com_out[1][46])
                                        );
                                        
                                        compress_module compress_303 (
                                            .x(u[1][47]),
                                            .d(10),
                                            .result(com_out[1][47])
                                        );
                                        
                                        compress_module compress_304 (
                                            .x(u[1][48]),
                                            .d(10),
                                            .result(com_out[1][48])
                                        );
                                        
                                        compress_module compress_305 (
                                            .x(u[1][49]),
                                            .d(10),
                                            .result(com_out[1][49])
                                        );
                                        
                                        compress_module compress_306 (
                                            .x(u[1][50]),
                                            .d(10),
                                            .result(com_out[1][50])
                                        );
                                        
                                        compress_module compress_307 (
                                            .x(u[1][51]),
                                            .d(10),
                                            .result(com_out[1][51])
                                        );
                                        
                                        compress_module compress_308 (
                                            .x(u[1][52]),
                                            .d(10),
                                            .result(com_out[1][52])
                                        );
                                        
                                        compress_module compress_309 (
                                            .x(u[1][53]),
                                            .d(10),
                                            .result(com_out[1][53])
                                        );
                                        
                                        compress_module compress_310 (
                                            .x(u[1][54]),
                                            .d(10),
                                            .result(com_out[1][54])
                                        );
                                        
                                        compress_module compress_311 (
                                            .x(u[1][55]),
                                            .d(10),
                                            .result(com_out[1][55])
                                        );
                                        
                                        compress_module compress_312 (
                                            .x(u[1][56]),
                                            .d(10),
                                            .result(com_out[1][56])
                                        );
                                        
                                        compress_module compress_313 (
                                            .x(u[1][57]),
                                            .d(10),
                                            .result(com_out[1][57])
                                        );
                                        
                                        compress_module compress_314 (
                                            .x(u[1][58]),
                                            .d(10),
                                            .result(com_out[1][58])
                                        );
                                        
                                        compress_module compress_315 (
                                            .x(u[1][59]),
                                            .d(10),
                                            .result(com_out[1][59])
                                        );
                                        
                                        compress_module compress_316 (
                                            .x(u[1][60]),
                                            .d(10),
                                            .result(com_out[1][60])
                                        );
                                        
                                        compress_module compress_317 (
                                            .x(u[1][61]),
                                            .d(10),
                                            .result(com_out[1][61])
                                        );
                                        
                                        compress_module compress_318 (
                                            .x(u[1][62]),
                                            .d(10),
                                            .result(com_out[1][62])
                                        );
                                        
                                        compress_module compress_319 (
                                            .x(u[1][63]),
                                            .d(10),
                                            .result(com_out[1][63])
                                        );
                                        
                                        compress_module compress_320 (
                                            .x(u[1][64]),
                                            .d(10),
                                            .result(com_out[1][64])
                                        );
                                        
                                        compress_module compress_321 (
                                            .x(u[1][65]),
                                            .d(10),
                                            .result(com_out[1][65])
                                        );
                                        
                                        compress_module compress_322 (
                                            .x(u[1][66]),
                                            .d(10),
                                            .result(com_out[1][66])
                                        );
                                        
                                        compress_module compress_323 (
                                            .x(u[1][67]),
                                            .d(10),
                                            .result(com_out[1][67])
                                        );
                                        
                                        compress_module compress_324 (
                                            .x(u[1][68]),
                                            .d(10),
                                            .result(com_out[1][68])
                                        );
                                        
                                        compress_module compress_325 (
                                            .x(u[1][69]),
                                            .d(10),
                                            .result(com_out[1][69])
                                        );
                                        
                                        compress_module compress_326 (
                                            .x(u[1][70]),
                                            .d(10),
                                            .result(com_out[1][70])
                                        );
                                        
                                        compress_module compress_327 (
                                            .x(u[1][71]),
                                            .d(10),
                                            .result(com_out[1][71])
                                        );
                                        
                                        compress_module compress_328 (
                                            .x(u[1][72]),
                                            .d(10),
                                            .result(com_out[1][72])
                                        );
                                        
                                        compress_module compress_329 (
                                            .x(u[1][73]),
                                            .d(10),
                                            .result(com_out[1][73])
                                        );
                                        
                                        compress_module compress_330 (
                                            .x(u[1][74]),
                                            .d(10),
                                            .result(com_out[1][74])
                                        );
                                        
                                        compress_module compress_331 (
                                            .x(u[1][75]),
                                            .d(10),
                                            .result(com_out[1][75])
                                        );
                                        
                                        compress_module compress_332 (
                                            .x(u[1][76]),
                                            .d(10),
                                            .result(com_out[1][76])
                                        );
                                        
                                        compress_module compress_333 (
                                            .x(u[1][77]),
                                            .d(10),
                                            .result(com_out[1][77])
                                        );
                                        
                                        compress_module compress_334 (
                                            .x(u[1][78]),
                                            .d(10),
                                            .result(com_out[1][78])
                                        );
                                        
                                        compress_module compress_335 (
                                            .x(u[1][79]),
                                            .d(10),
                                            .result(com_out[1][79])
                                        );
                                        
                                        compress_module compress_336 (
                                            .x(u[1][80]),
                                            .d(10),
                                            .result(com_out[1][80])
                                        );
                                        
                                        compress_module compress_337 (
                                            .x(u[1][81]),
                                            .d(10),
                                            .result(com_out[1][81])
                                        );
                                        
                                        compress_module compress_338 (
                                            .x(u[1][82]),
                                            .d(10),
                                            .result(com_out[1][82])
                                        );
                                        
                                        compress_module compress_339 (
                                            .x(u[1][83]),
                                            .d(10),
                                            .result(com_out[1][83])
                                        );
                                        
                                        compress_module compress_340 (
                                            .x(u[1][84]),
                                            .d(10),
                                            .result(com_out[1][84])
                                        );
                                        
                                        compress_module compress_341 (
                                            .x(u[1][85]),
                                            .d(10),
                                            .result(com_out[1][85])
                                        );
                                        
                                        compress_module compress_342 (
                                            .x(u[1][86]),
                                            .d(10),
                                            .result(com_out[1][86])
                                        );
                                        
                                        compress_module compress_343 (
                                            .x(u[1][87]),
                                            .d(10),
                                            .result(com_out[1][87])
                                        );
                                        
                                        compress_module compress_344 (
                                            .x(u[1][88]),
                                            .d(10),
                                            .result(com_out[1][88])
                                        );
                                        
                                        compress_module compress_345 (
                                            .x(u[1][89]),
                                            .d(10),
                                            .result(com_out[1][89])
                                        );
                                        
                                        compress_module compress_346 (
                                            .x(u[1][90]),
                                            .d(10),
                                            .result(com_out[1][90])
                                        );
                                        
                                        compress_module compress_347 (
                                            .x(u[1][91]),
                                            .d(10),
                                            .result(com_out[1][91])
                                        );
                                        
                                        compress_module compress_348 (
                                            .x(u[1][92]),
                                            .d(10),
                                            .result(com_out[1][92])
                                        );
                                        
                                        compress_module compress_349 (
                                            .x(u[1][93]),
                                            .d(10),
                                            .result(com_out[1][93])
                                        );
                                        
                                        compress_module compress_350 (
                                            .x(u[1][94]),
                                            .d(10),
                                            .result(com_out[1][94])
                                        );
                                        
                                        compress_module compress_351 (
                                            .x(u[1][95]),
                                            .d(10),
                                            .result(com_out[1][95])
                                        );
                                        
                                        compress_module compress_352 (
                                            .x(u[1][96]),
                                            .d(10),
                                            .result(com_out[1][96])
                                        );
                                        
                                        compress_module compress_353 (
                                            .x(u[1][97]),
                                            .d(10),
                                            .result(com_out[1][97])
                                        );
                                        
                                        compress_module compress_354 (
                                            .x(u[1][98]),
                                            .d(10),
                                            .result(com_out[1][98])
                                        );
                                        
                                        compress_module compress_355 (
                                            .x(u[1][99]),
                                            .d(10),
                                            .result(com_out[1][99])
                                        );
                                        
                                        compress_module compress_356 (
                                            .x(u[1][100]),
                                            .d(10),
                                            .result(com_out[1][100])
                                        );
                                        
                                        compress_module compress_357 (
                                            .x(u[1][101]),
                                            .d(10),
                                            .result(com_out[1][101])
                                        );
                                        
                                        compress_module compress_358 (
                                            .x(u[1][102]),
                                            .d(10),
                                            .result(com_out[1][102])
                                        );
                                        
                                        compress_module compress_359 (
                                            .x(u[1][103]),
                                            .d(10),
                                            .result(com_out[1][103])
                                        );
                                        
                                        compress_module compress_360 (
                                            .x(u[1][104]),
                                            .d(10),
                                            .result(com_out[1][104])
                                        );
                                        
                                        compress_module compress_361 (
                                            .x(u[1][105]),
                                            .d(10),
                                            .result(com_out[1][105])
                                        );
                                        
                                        compress_module compress_362 (
                                            .x(u[1][106]),
                                            .d(10),
                                            .result(com_out[1][106])
                                        );
                                        
                                        compress_module compress_363 (
                                            .x(u[1][107]),
                                            .d(10),
                                            .result(com_out[1][107])
                                        );
                                        
                                        compress_module compress_364 (
                                            .x(u[1][108]),
                                            .d(10),
                                            .result(com_out[1][108])
                                        );
                                        
                                        compress_module compress_365 (
                                            .x(u[1][109]),
                                            .d(10),
                                            .result(com_out[1][109])
                                        );
                                        
                                        compress_module compress_366 (
                                            .x(u[1][110]),
                                            .d(10),
                                            .result(com_out[1][110])
                                        );
                                        
                                        compress_module compress_367 (
                                            .x(u[1][111]),
                                            .d(10),
                                            .result(com_out[1][111])
                                        );
                                        
                                        compress_module compress_368 (
                                            .x(u[1][112]),
                                            .d(10),
                                            .result(com_out[1][112])
                                        );
                                        
                                        compress_module compress_369 (
                                            .x(u[1][113]),
                                            .d(10),
                                            .result(com_out[1][113])
                                        );
                                        
                                        compress_module compress_370 (
                                            .x(u[1][114]),
                                            .d(10),
                                            .result(com_out[1][114])
                                        );
                                        
                                        compress_module compress_371 (
                                            .x(u[1][115]),
                                            .d(10),
                                            .result(com_out[1][115])
                                        );
                                        
                                        compress_module compress_372 (
                                            .x(u[1][116]),
                                            .d(10),
                                            .result(com_out[1][116])
                                        );
                                        
                                        compress_module compress_373 (
                                            .x(u[1][117]),
                                            .d(10),
                                            .result(com_out[1][117])
                                        );
                                        
                                        compress_module compress_374 (
                                            .x(u[1][118]),
                                            .d(10),
                                            .result(com_out[1][118])
                                        );
                                        
                                        compress_module compress_375 (
                                            .x(u[1][119]),
                                            .d(10),
                                            .result(com_out[1][119])
                                        );
                                        
                                        compress_module compress_376 (
                                            .x(u[1][120]),
                                            .d(10),
                                            .result(com_out[1][120])
                                        );
                                        
                                        compress_module compress_377 (
                                            .x(u[1][121]),
                                            .d(10),
                                            .result(com_out[1][121])
                                        );
                                        
                                        compress_module compress_378 (
                                            .x(u[1][122]),
                                            .d(10),
                                            .result(com_out[1][122])
                                        );
                                        
                                        compress_module compress_379 (
                                            .x(u[1][123]),
                                            .d(10),
                                            .result(com_out[1][123])
                                        );
                                        
                                        compress_module compress_380 (
                                            .x(u[1][124]),
                                            .d(10),
                                            .result(com_out[1][124])
                                        );
                                        
                                        compress_module compress_381 (
                                            .x(u[1][125]),
                                            .d(10),
                                            .result(com_out[1][125])
                                        );
                                        
                                        compress_module compress_382 (
                                            .x(u[1][126]),
                                            .d(10),
                                            .result(com_out[1][126])
                                        );
                                        
                                        compress_module compress_383 (
                                            .x(u[1][127]),
                                            .d(10),
                                            .result(com_out[1][127])
                                        );
                                        
                                        compress_module compress_384 (
                                            .x(u[1][128]),
                                            .d(10),
                                            .result(com_out[1][128])
                                        );
                                        
                                        compress_module compress_385 (
                                            .x(u[1][129]),
                                            .d(10),
                                            .result(com_out[1][129])
                                        );
                                        
                                        compress_module compress_386 (
                                            .x(u[1][130]),
                                            .d(10),
                                            .result(com_out[1][130])
                                        );
                                        
                                        compress_module compress_387 (
                                            .x(u[1][131]),
                                            .d(10),
                                            .result(com_out[1][131])
                                        );
                                        
                                        compress_module compress_388 (
                                            .x(u[1][132]),
                                            .d(10),
                                            .result(com_out[1][132])
                                        );
                                        
                                        compress_module compress_389 (
                                            .x(u[1][133]),
                                            .d(10),
                                            .result(com_out[1][133])
                                        );
                                        
                                        compress_module compress_390 (
                                            .x(u[1][134]),
                                            .d(10),
                                            .result(com_out[1][134])
                                        );
                                        
                                        compress_module compress_391 (
                                            .x(u[1][135]),
                                            .d(10),
                                            .result(com_out[1][135])
                                        );
                                        
                                        compress_module compress_392 (
                                            .x(u[1][136]),
                                            .d(10),
                                            .result(com_out[1][136])
                                        );
                                        
                                        compress_module compress_393 (
                                            .x(u[1][137]),
                                            .d(10),
                                            .result(com_out[1][137])
                                        );
                                        
                                        compress_module compress_394 (
                                            .x(u[1][138]),
                                            .d(10),
                                            .result(com_out[1][138])
                                        );
                                        
                                        compress_module compress_395 (
                                            .x(u[1][139]),
                                            .d(10),
                                            .result(com_out[1][139])
                                        );
                                        
                                        compress_module compress_396 (
                                            .x(u[1][140]),
                                            .d(10),
                                            .result(com_out[1][140])
                                        );
                                        
                                        compress_module compress_397 (
                                            .x(u[1][141]),
                                            .d(10),
                                            .result(com_out[1][141])
                                        );
                                        
                                        compress_module compress_398 (
                                            .x(u[1][142]),
                                            .d(10),
                                            .result(com_out[1][142])
                                        );
                                        
                                        compress_module compress_399 (
                                            .x(u[1][143]),
                                            .d(10),
                                            .result(com_out[1][143])
                                        );
                                        
                                        compress_module compress_400 (
                                            .x(u[1][144]),
                                            .d(10),
                                            .result(com_out[1][144])
                                        );
                                        
                                        compress_module compress_401 (
                                            .x(u[1][145]),
                                            .d(10),
                                            .result(com_out[1][145])
                                        );
                                        
                                        compress_module compress_402 (
                                            .x(u[1][146]),
                                            .d(10),
                                            .result(com_out[1][146])
                                        );
                                        
                                        compress_module compress_403 (
                                            .x(u[1][147]),
                                            .d(10),
                                            .result(com_out[1][147])
                                        );
                                        
                                        compress_module compress_404 (
                                            .x(u[1][148]),
                                            .d(10),
                                            .result(com_out[1][148])
                                        );
                                        
                                        compress_module compress_405 (
                                            .x(u[1][149]),
                                            .d(10),
                                            .result(com_out[1][149])
                                        );
                                        
                                        compress_module compress_406 (
                                            .x(u[1][150]),
                                            .d(10),
                                            .result(com_out[1][150])
                                        );
                                        
                                        compress_module compress_407 (
                                            .x(u[1][151]),
                                            .d(10),
                                            .result(com_out[1][151])
                                        );
                                        
                                        compress_module compress_408 (
                                            .x(u[1][152]),
                                            .d(10),
                                            .result(com_out[1][152])
                                        );
                                        
                                        compress_module compress_409 (
                                            .x(u[1][153]),
                                            .d(10),
                                            .result(com_out[1][153])
                                        );
                                        
                                        compress_module compress_410 (
                                            .x(u[1][154]),
                                            .d(10),
                                            .result(com_out[1][154])
                                        );
                                        
                                        compress_module compress_411 (
                                            .x(u[1][155]),
                                            .d(10),
                                            .result(com_out[1][155])
                                        );
                                        
                                        compress_module compress_412 (
                                            .x(u[1][156]),
                                            .d(10),
                                            .result(com_out[1][156])
                                        );
                                        
                                        compress_module compress_413 (
                                            .x(u[1][157]),
                                            .d(10),
                                            .result(com_out[1][157])
                                        );
                                        
                                        compress_module compress_414 (
                                            .x(u[1][158]),
                                            .d(10),
                                            .result(com_out[1][158])
                                        );
                                        
                                        compress_module compress_415 (
                                            .x(u[1][159]),
                                            .d(10),
                                            .result(com_out[1][159])
                                        );
                                        
                                        compress_module compress_416 (
                                            .x(u[1][160]),
                                            .d(10),
                                            .result(com_out[1][160])
                                        );
                                        
                                        compress_module compress_417 (
                                            .x(u[1][161]),
                                            .d(10),
                                            .result(com_out[1][161])
                                        );
                                        
                                        compress_module compress_418 (
                                            .x(u[1][162]),
                                            .d(10),
                                            .result(com_out[1][162])
                                        );
                                        
                                        compress_module compress_419 (
                                            .x(u[1][163]),
                                            .d(10),
                                            .result(com_out[1][163])
                                        );
                                        
                                        compress_module compress_420 (
                                            .x(u[1][164]),
                                            .d(10),
                                            .result(com_out[1][164])
                                        );
                                        
                                        compress_module compress_421 (
                                            .x(u[1][165]),
                                            .d(10),
                                            .result(com_out[1][165])
                                        );
                                        
                                        compress_module compress_422 (
                                            .x(u[1][166]),
                                            .d(10),
                                            .result(com_out[1][166])
                                        );
                                        
                                        compress_module compress_423 (
                                            .x(u[1][167]),
                                            .d(10),
                                            .result(com_out[1][167])
                                        );
                                        
                                        compress_module compress_424 (
                                            .x(u[1][168]),
                                            .d(10),
                                            .result(com_out[1][168])
                                        );
                                        
                                        compress_module compress_425 (
                                            .x(u[1][169]),
                                            .d(10),
                                            .result(com_out[1][169])
                                        );
                                        
                                        compress_module compress_426 (
                                            .x(u[1][170]),
                                            .d(10),
                                            .result(com_out[1][170])
                                        );
                                        
                                        compress_module compress_427 (
                                            .x(u[1][171]),
                                            .d(10),
                                            .result(com_out[1][171])
                                        );
                                        
                                        compress_module compress_428 (
                                            .x(u[1][172]),
                                            .d(10),
                                            .result(com_out[1][172])
                                        );
                                        
                                        compress_module compress_429 (
                                            .x(u[1][173]),
                                            .d(10),
                                            .result(com_out[1][173])
                                        );
                                        
                                        compress_module compress_430 (
                                            .x(u[1][174]),
                                            .d(10),
                                            .result(com_out[1][174])
                                        );
                                        
                                        compress_module compress_431 (
                                            .x(u[1][175]),
                                            .d(10),
                                            .result(com_out[1][175])
                                        );
                                        
                                        compress_module compress_432 (
                                            .x(u[1][176]),
                                            .d(10),
                                            .result(com_out[1][176])
                                        );
                                        
                                        compress_module compress_433 (
                                            .x(u[1][177]),
                                            .d(10),
                                            .result(com_out[1][177])
                                        );
                                        
                                        compress_module compress_434 (
                                            .x(u[1][178]),
                                            .d(10),
                                            .result(com_out[1][178])
                                        );
                                        
                                        compress_module compress_435 (
                                            .x(u[1][179]),
                                            .d(10),
                                            .result(com_out[1][179])
                                        );
                                        
                                        compress_module compress_436 (
                                            .x(u[1][180]),
                                            .d(10),
                                            .result(com_out[1][180])
                                        );
                                        
                                        compress_module compress_437 (
                                            .x(u[1][181]),
                                            .d(10),
                                            .result(com_out[1][181])
                                        );
                                        
                                        compress_module compress_438 (
                                            .x(u[1][182]),
                                            .d(10),
                                            .result(com_out[1][182])
                                        );
                                        
                                        compress_module compress_439 (
                                            .x(u[1][183]),
                                            .d(10),
                                            .result(com_out[1][183])
                                        );
                                        
                                        compress_module compress_440 (
                                            .x(u[1][184]),
                                            .d(10),
                                            .result(com_out[1][184])
                                        );
                                        
                                        compress_module compress_441 (
                                            .x(u[1][185]),
                                            .d(10),
                                            .result(com_out[1][185])
                                        );
                                        
                                        compress_module compress_442 (
                                            .x(u[1][186]),
                                            .d(10),
                                            .result(com_out[1][186])
                                        );
                                        
                                        compress_module compress_443 (
                                            .x(u[1][187]),
                                            .d(10),
                                            .result(com_out[1][187])
                                        );
                                        
                                        compress_module compress_444 (
                                            .x(u[1][188]),
                                            .d(10),
                                            .result(com_out[1][188])
                                        );
                                        
                                        compress_module compress_445 (
                                            .x(u[1][189]),
                                            .d(10),
                                            .result(com_out[1][189])
                                        );
                                        
                                        compress_module compress_446 (
                                            .x(u[1][190]),
                                            .d(10),
                                            .result(com_out[1][190])
                                        );
                                        
                                        compress_module compress_447 (
                                            .x(u[1][191]),
                                            .d(10),
                                            .result(com_out[1][191])
                                        );
                                        
                                        compress_module compress_448 (
                                            .x(u[1][192]),
                                            .d(10),
                                            .result(com_out[1][192])
                                        );
                                        
                                        compress_module compress_449 (
                                            .x(u[1][193]),
                                            .d(10),
                                            .result(com_out[1][193])
                                        );
                                        
                                        compress_module compress_450 (
                                            .x(u[1][194]),
                                            .d(10),
                                            .result(com_out[1][194])
                                        );
                                        
                                        compress_module compress_451 (
                                            .x(u[1][195]),
                                            .d(10),
                                            .result(com_out[1][195])
                                        );
                                        
                                        compress_module compress_452 (
                                            .x(u[1][196]),
                                            .d(10),
                                            .result(com_out[1][196])
                                        );
                                        
                                        compress_module compress_453 (
                                            .x(u[1][197]),
                                            .d(10),
                                            .result(com_out[1][197])
                                        );
                                        
                                        compress_module compress_454 (
                                            .x(u[1][198]),
                                            .d(10),
                                            .result(com_out[1][198])
                                        );
                                        
                                        compress_module compress_455 (
                                            .x(u[1][199]),
                                            .d(10),
                                            .result(com_out[1][199])
                                        );
                                        
                                        compress_module compress_456 (
                                            .x(u[1][200]),
                                            .d(10),
                                            .result(com_out[1][200])
                                        );
                                        
                                        compress_module compress_457 (
                                            .x(u[1][201]),
                                            .d(10),
                                            .result(com_out[1][201])
                                        );
                                        
                                        compress_module compress_458 (
                                            .x(u[1][202]),
                                            .d(10),
                                            .result(com_out[1][202])
                                        );
                                        
                                        compress_module compress_459 (
                                            .x(u[1][203]),
                                            .d(10),
                                            .result(com_out[1][203])
                                        );
                                        
                                        compress_module compress_460 (
                                            .x(u[1][204]),
                                            .d(10),
                                            .result(com_out[1][204])
                                        );
                                        
                                        compress_module compress_461 (
                                            .x(u[1][205]),
                                            .d(10),
                                            .result(com_out[1][205])
                                        );
                                        
                                        compress_module compress_462 (
                                            .x(u[1][206]),
                                            .d(10),
                                            .result(com_out[1][206])
                                        );
                                        
                                        compress_module compress_463 (
                                            .x(u[1][207]),
                                            .d(10),
                                            .result(com_out[1][207])
                                        );
                                        
                                        compress_module compress_464 (
                                            .x(u[1][208]),
                                            .d(10),
                                            .result(com_out[1][208])
                                        );
                                        
                                        compress_module compress_465 (
                                            .x(u[1][209]),
                                            .d(10),
                                            .result(com_out[1][209])
                                        );
                                        
                                        compress_module compress_466 (
                                            .x(u[1][210]),
                                            .d(10),
                                            .result(com_out[1][210])
                                        );
                                        
                                        compress_module compress_467 (
                                            .x(u[1][211]),
                                            .d(10),
                                            .result(com_out[1][211])
                                        );
                                        
                                        compress_module compress_468 (
                                            .x(u[1][212]),
                                            .d(10),
                                            .result(com_out[1][212])
                                        );
                                        
                                        compress_module compress_469 (
                                            .x(u[1][213]),
                                            .d(10),
                                            .result(com_out[1][213])
                                        );
                                        
                                        compress_module compress_470 (
                                            .x(u[1][214]),
                                            .d(10),
                                            .result(com_out[1][214])
                                        );
                                        
                                        compress_module compress_471 (
                                            .x(u[1][215]),
                                            .d(10),
                                            .result(com_out[1][215])
                                        );
                                        
                                        compress_module compress_472 (
                                            .x(u[1][216]),
                                            .d(10),
                                            .result(com_out[1][216])
                                        );
                                        
                                        compress_module compress_473 (
                                            .x(u[1][217]),
                                            .d(10),
                                            .result(com_out[1][217])
                                        );
                                        
                                        compress_module compress_474 (
                                            .x(u[1][218]),
                                            .d(10),
                                            .result(com_out[1][218])
                                        );
                                        
                                        compress_module compress_475 (
                                            .x(u[1][219]),
                                            .d(10),
                                            .result(com_out[1][219])
                                        );
                                        
                                        compress_module compress_476 (
                                            .x(u[1][220]),
                                            .d(10),
                                            .result(com_out[1][220])
                                        );
                                        
                                        compress_module compress_477 (
                                            .x(u[1][221]),
                                            .d(10),
                                            .result(com_out[1][221])
                                        );
                                        
                                        compress_module compress_478 (
                                            .x(u[1][222]),
                                            .d(10),
                                            .result(com_out[1][222])
                                        );
                                        
                                        compress_module compress_479 (
                                            .x(u[1][223]),
                                            .d(10),
                                            .result(com_out[1][223])
                                        );
                                        
                                        compress_module compress_480 (
                                            .x(u[1][224]),
                                            .d(10),
                                            .result(com_out[1][224])
                                        );
                                        
                                        compress_module compress_481 (
                                            .x(u[1][225]),
                                            .d(10),
                                            .result(com_out[1][225])
                                        );
                                        
                                        compress_module compress_482 (
                                            .x(u[1][226]),
                                            .d(10),
                                            .result(com_out[1][226])
                                        );
                                        
                                        compress_module compress_483 (
                                            .x(u[1][227]),
                                            .d(10),
                                            .result(com_out[1][227])
                                        );
                                        
                                        compress_module compress_484 (
                                            .x(u[1][228]),
                                            .d(10),
                                            .result(com_out[1][228])
                                        );
                                        
                                        compress_module compress_485 (
                                            .x(u[1][229]),
                                            .d(10),
                                            .result(com_out[1][229])
                                        );
                                        
                                        compress_module compress_486 (
                                            .x(u[1][230]),
                                            .d(10),
                                            .result(com_out[1][230])
                                        );
                                        
                                        compress_module compress_487 (
                                            .x(u[1][231]),
                                            .d(10),
                                            .result(com_out[1][231])
                                        );
                                        
                                        compress_module compress_488 (
                                            .x(u[1][232]),
                                            .d(10),
                                            .result(com_out[1][232])
                                        );
                                        
                                        compress_module compress_489 (
                                            .x(u[1][233]),
                                            .d(10),
                                            .result(com_out[1][233])
                                        );
                                        
                                        compress_module compress_490 (
                                            .x(u[1][234]),
                                            .d(10),
                                            .result(com_out[1][234])
                                        );
                                        
                                        compress_module compress_491 (
                                            .x(u[1][235]),
                                            .d(10),
                                            .result(com_out[1][235])
                                        );
                                        
                                        compress_module compress_492 (
                                            .x(u[1][236]),
                                            .d(10),
                                            .result(com_out[1][236])
                                        );
                                        
                                        compress_module compress_493 (
                                            .x(u[1][237]),
                                            .d(10),
                                            .result(com_out[1][237])
                                        );
                                        
                                        compress_module compress_494 (
                                            .x(u[1][238]),
                                            .d(10),
                                            .result(com_out[1][238])
                                        );
                                        
                                        compress_module compress_495 (
                                            .x(u[1][239]),
                                            .d(10),
                                            .result(com_out[1][239])
                                        );
                                        
                                        compress_module compress_496 (
                                            .x(u[1][240]),
                                            .d(10),
                                            .result(com_out[1][240])
                                        );
                                        
                                        compress_module compress_497 (
                                            .x(u[1][241]),
                                            .d(10),
                                            .result(com_out[1][241])
                                        );
                                        
                                        compress_module compress_498 (
                                            .x(u[1][242]),
                                            .d(10),
                                            .result(com_out[1][242])
                                        );
                                        
                                        compress_module compress_499 (
                                            .x(u[1][243]),
                                            .d(10),
                                            .result(com_out[1][243])
                                        );
                                        
                                        compress_module compress_500 (
                                            .x(u[1][244]),
                                            .d(10),
                                            .result(com_out[1][244])
                                        );
                                        
                                        compress_module compress_501 (
                                            .x(u[1][245]),
                                            .d(10),
                                            .result(com_out[1][245])
                                        );
                                        
                                        compress_module compress_502 (
                                            .x(u[1][246]),
                                            .d(10),
                                            .result(com_out[1][246])
                                        );
                                        
                                        compress_module compress_503 (
                                            .x(u[1][247]),
                                            .d(10),
                                            .result(com_out[1][247])
                                        );
                                        
                                        compress_module compress_504 (
                                            .x(u[1][248]),
                                            .d(10),
                                            .result(com_out[1][248])
                                        );
                                        
                                        compress_module compress_505 (
                                            .x(u[1][249]),
                                            .d(10),
                                            .result(com_out[1][249])
                                        );
                                        
                                        compress_module compress_506 (
                                            .x(u[1][250]),
                                            .d(10),
                                            .result(com_out[1][250])
                                        );
                                        
                                        compress_module compress_507 (
                                            .x(u[1][251]),
                                            .d(10),
                                            .result(com_out[1][251])
                                        );
                                        
                                        compress_module compress_508 (
                                            .x(u[1][252]),
                                            .d(10),
                                            .result(com_out[1][252])
                                        );
                                        
                                        compress_module compress_509 (
                                            .x(u[1][253]),
                                            .d(10),
                                            .result(com_out[1][253])
                                        );
                                        
                                        compress_module compress_510 (
                                            .x(u[1][254]),
                                            .d(10),
                                            .result(com_out[1][254])
                                        );
                                        
                                        compress_module compress_511 (
                                            .x(u[1][255]),
                                            .d(10),
                                            .result(com_out[1][255])
                                        );
                                        
                                        compress_module compress_512 (
                                            .x(u[2][0]),
                                            .d(10),
                                            .result(com_out[2][0])
                                        );
                                        
                                        compress_module compress_513 (
                                            .x(u[2][1]),
                                            .d(10),
                                            .result(com_out[2][1])
                                        );
                                        
                                        compress_module compress_514 (
                                            .x(u[2][2]),
                                            .d(10),
                                            .result(com_out[2][2])
                                        );
                                        
                                        compress_module compress_515 (
                                            .x(u[2][3]),
                                            .d(10),
                                            .result(com_out[2][3])
                                        );
                                        
                                        compress_module compress_516 (
                                            .x(u[2][4]),
                                            .d(10),
                                            .result(com_out[2][4])
                                        );
                                        
                                        compress_module compress_517 (
                                            .x(u[2][5]),
                                            .d(10),
                                            .result(com_out[2][5])
                                        );
                                        
                                        compress_module compress_518 (
                                            .x(u[2][6]),
                                            .d(10),
                                            .result(com_out[2][6])
                                        );
                                        
                                        compress_module compress_519 (
                                            .x(u[2][7]),
                                            .d(10),
                                            .result(com_out[2][7])
                                        );
                                        
                                        compress_module compress_520 (
                                            .x(u[2][8]),
                                            .d(10),
                                            .result(com_out[2][8])
                                        );
                                        
                                        compress_module compress_521 (
                                            .x(u[2][9]),
                                            .d(10),
                                            .result(com_out[2][9])
                                        );
                                        
                                        compress_module compress_522 (
                                            .x(u[2][10]),
                                            .d(10),
                                            .result(com_out[2][10])
                                        );
                                        
                                        compress_module compress_523 (
                                            .x(u[2][11]),
                                            .d(10),
                                            .result(com_out[2][11])
                                        );
                                        
                                        compress_module compress_524 (
                                            .x(u[2][12]),
                                            .d(10),
                                            .result(com_out[2][12])
                                        );
                                        
                                        compress_module compress_525 (
                                            .x(u[2][13]),
                                            .d(10),
                                            .result(com_out[2][13])
                                        );
                                        
                                        compress_module compress_526 (
                                            .x(u[2][14]),
                                            .d(10),
                                            .result(com_out[2][14])
                                        );
                                        
                                        compress_module compress_527 (
                                            .x(u[2][15]),
                                            .d(10),
                                            .result(com_out[2][15])
                                        );
                                        
                                        compress_module compress_528 (
                                            .x(u[2][16]),
                                            .d(10),
                                            .result(com_out[2][16])
                                        );
                                        
                                        compress_module compress_529 (
                                            .x(u[2][17]),
                                            .d(10),
                                            .result(com_out[2][17])
                                        );
                                        
                                        compress_module compress_530 (
                                            .x(u[2][18]),
                                            .d(10),
                                            .result(com_out[2][18])
                                        );
                                        
                                        compress_module compress_531 (
                                            .x(u[2][19]),
                                            .d(10),
                                            .result(com_out[2][19])
                                        );
                                        
                                        compress_module compress_532 (
                                            .x(u[2][20]),
                                            .d(10),
                                            .result(com_out[2][20])
                                        );
                                        
                                        compress_module compress_533 (
                                            .x(u[2][21]),
                                            .d(10),
                                            .result(com_out[2][21])
                                        );
                                        
                                        compress_module compress_534 (
                                            .x(u[2][22]),
                                            .d(10),
                                            .result(com_out[2][22])
                                        );
                                        
                                        compress_module compress_535 (
                                            .x(u[2][23]),
                                            .d(10),
                                            .result(com_out[2][23])
                                        );
                                        
                                        compress_module compress_536 (
                                            .x(u[2][24]),
                                            .d(10),
                                            .result(com_out[2][24])
                                        );
                                        
                                        compress_module compress_537 (
                                            .x(u[2][25]),
                                            .d(10),
                                            .result(com_out[2][25])
                                        );
                                        
                                        compress_module compress_538 (
                                            .x(u[2][26]),
                                            .d(10),
                                            .result(com_out[2][26])
                                        );
                                        
                                        compress_module compress_539 (
                                            .x(u[2][27]),
                                            .d(10),
                                            .result(com_out[2][27])
                                        );
                                        
                                        compress_module compress_540 (
                                            .x(u[2][28]),
                                            .d(10),
                                            .result(com_out[2][28])
                                        );
                                        
                                        compress_module compress_541 (
                                            .x(u[2][29]),
                                            .d(10),
                                            .result(com_out[2][29])
                                        );
                                        
                                        compress_module compress_542 (
                                            .x(u[2][30]),
                                            .d(10),
                                            .result(com_out[2][30])
                                        );
                                        
                                        compress_module compress_543 (
                                            .x(u[2][31]),
                                            .d(10),
                                            .result(com_out[2][31])
                                        );
                                        
                                        compress_module compress_544 (
                                            .x(u[2][32]),
                                            .d(10),
                                            .result(com_out[2][32])
                                        );
                                        
                                        compress_module compress_545 (
                                            .x(u[2][33]),
                                            .d(10),
                                            .result(com_out[2][33])
                                        );
                                        
                                        compress_module compress_546 (
                                            .x(u[2][34]),
                                            .d(10),
                                            .result(com_out[2][34])
                                        );
                                        
                                        compress_module compress_547 (
                                            .x(u[2][35]),
                                            .d(10),
                                            .result(com_out[2][35])
                                        );
                                        
                                        compress_module compress_548 (
                                            .x(u[2][36]),
                                            .d(10),
                                            .result(com_out[2][36])
                                        );
                                        
                                        compress_module compress_549 (
                                            .x(u[2][37]),
                                            .d(10),
                                            .result(com_out[2][37])
                                        );
                                        
                                        compress_module compress_550 (
                                            .x(u[2][38]),
                                            .d(10),
                                            .result(com_out[2][38])
                                        );
                                        
                                        compress_module compress_551 (
                                            .x(u[2][39]),
                                            .d(10),
                                            .result(com_out[2][39])
                                        );
                                        
                                        compress_module compress_552 (
                                            .x(u[2][40]),
                                            .d(10),
                                            .result(com_out[2][40])
                                        );
                                        
                                        compress_module compress_553 (
                                            .x(u[2][41]),
                                            .d(10),
                                            .result(com_out[2][41])
                                        );
                                        
                                        compress_module compress_554 (
                                            .x(u[2][42]),
                                            .d(10),
                                            .result(com_out[2][42])
                                        );
                                        
                                        compress_module compress_555 (
                                            .x(u[2][43]),
                                            .d(10),
                                            .result(com_out[2][43])
                                        );
                                        
                                        compress_module compress_556 (
                                            .x(u[2][44]),
                                            .d(10),
                                            .result(com_out[2][44])
                                        );
                                        
                                        compress_module compress_557 (
                                            .x(u[2][45]),
                                            .d(10),
                                            .result(com_out[2][45])
                                        );
                                        
                                        compress_module compress_558 (
                                            .x(u[2][46]),
                                            .d(10),
                                            .result(com_out[2][46])
                                        );
                                        
                                        compress_module compress_559 (
                                            .x(u[2][47]),
                                            .d(10),
                                            .result(com_out[2][47])
                                        );
                                        
                                        compress_module compress_560 (
                                            .x(u[2][48]),
                                            .d(10),
                                            .result(com_out[2][48])
                                        );
                                        
                                        compress_module compress_561 (
                                            .x(u[2][49]),
                                            .d(10),
                                            .result(com_out[2][49])
                                        );
                                        
                                        compress_module compress_562 (
                                            .x(u[2][50]),
                                            .d(10),
                                            .result(com_out[2][50])
                                        );
                                        
                                        compress_module compress_563 (
                                            .x(u[2][51]),
                                            .d(10),
                                            .result(com_out[2][51])
                                        );
                                        
                                        compress_module compress_564 (
                                            .x(u[2][52]),
                                            .d(10),
                                            .result(com_out[2][52])
                                        );
                                        
                                        compress_module compress_565 (
                                            .x(u[2][53]),
                                            .d(10),
                                            .result(com_out[2][53])
                                        );
                                        
                                        compress_module compress_566 (
                                            .x(u[2][54]),
                                            .d(10),
                                            .result(com_out[2][54])
                                        );
                                        
                                        compress_module compress_567 (
                                            .x(u[2][55]),
                                            .d(10),
                                            .result(com_out[2][55])
                                        );
                                        
                                        compress_module compress_568 (
                                            .x(u[2][56]),
                                            .d(10),
                                            .result(com_out[2][56])
                                        );
                                        
                                        compress_module compress_569 (
                                            .x(u[2][57]),
                                            .d(10),
                                            .result(com_out[2][57])
                                        );
                                        
                                        compress_module compress_570 (
                                            .x(u[2][58]),
                                            .d(10),
                                            .result(com_out[2][58])
                                        );
                                        
                                        compress_module compress_571 (
                                            .x(u[2][59]),
                                            .d(10),
                                            .result(com_out[2][59])
                                        );
                                        
                                        compress_module compress_572 (
                                            .x(u[2][60]),
                                            .d(10),
                                            .result(com_out[2][60])
                                        );
                                        
                                        compress_module compress_573 (
                                            .x(u[2][61]),
                                            .d(10),
                                            .result(com_out[2][61])
                                        );
                                        
                                        compress_module compress_574 (
                                            .x(u[2][62]),
                                            .d(10),
                                            .result(com_out[2][62])
                                        );
                                        
                                        compress_module compress_575 (
                                            .x(u[2][63]),
                                            .d(10),
                                            .result(com_out[2][63])
                                        );
                                        
                                        compress_module compress_576 (
                                            .x(u[2][64]),
                                            .d(10),
                                            .result(com_out[2][64])
                                        );
                                        
                                        compress_module compress_577 (
                                            .x(u[2][65]),
                                            .d(10),
                                            .result(com_out[2][65])
                                        );
                                        
                                        compress_module compress_578 (
                                            .x(u[2][66]),
                                            .d(10),
                                            .result(com_out[2][66])
                                        );
                                        
                                        compress_module compress_579 (
                                            .x(u[2][67]),
                                            .d(10),
                                            .result(com_out[2][67])
                                        );
                                        
                                        compress_module compress_580 (
                                            .x(u[2][68]),
                                            .d(10),
                                            .result(com_out[2][68])
                                        );
                                        
                                        compress_module compress_581 (
                                            .x(u[2][69]),
                                            .d(10),
                                            .result(com_out[2][69])
                                        );
                                        
                                        compress_module compress_582 (
                                            .x(u[2][70]),
                                            .d(10),
                                            .result(com_out[2][70])
                                        );
                                        
                                        compress_module compress_583 (
                                            .x(u[2][71]),
                                            .d(10),
                                            .result(com_out[2][71])
                                        );
                                        
                                        compress_module compress_584 (
                                            .x(u[2][72]),
                                            .d(10),
                                            .result(com_out[2][72])
                                        );
                                        
                                        compress_module compress_585 (
                                            .x(u[2][73]),
                                            .d(10),
                                            .result(com_out[2][73])
                                        );
                                        
                                        compress_module compress_586 (
                                            .x(u[2][74]),
                                            .d(10),
                                            .result(com_out[2][74])
                                        );
                                        
                                        compress_module compress_587 (
                                            .x(u[2][75]),
                                            .d(10),
                                            .result(com_out[2][75])
                                        );
                                        
                                        compress_module compress_588 (
                                            .x(u[2][76]),
                                            .d(10),
                                            .result(com_out[2][76])
                                        );
                                        
                                        compress_module compress_589 (
                                            .x(u[2][77]),
                                            .d(10),
                                            .result(com_out[2][77])
                                        );
                                        
                                        compress_module compress_590 (
                                            .x(u[2][78]),
                                            .d(10),
                                            .result(com_out[2][78])
                                        );
                                        
                                        compress_module compress_591 (
                                            .x(u[2][79]),
                                            .d(10),
                                            .result(com_out[2][79])
                                        );
                                        
                                        compress_module compress_592 (
                                            .x(u[2][80]),
                                            .d(10),
                                            .result(com_out[2][80])
                                        );
                                        
                                        compress_module compress_593 (
                                            .x(u[2][81]),
                                            .d(10),
                                            .result(com_out[2][81])
                                        );
                                        
                                        compress_module compress_594 (
                                            .x(u[2][82]),
                                            .d(10),
                                            .result(com_out[2][82])
                                        );
                                        
                                        compress_module compress_595 (
                                            .x(u[2][83]),
                                            .d(10),
                                            .result(com_out[2][83])
                                        );
                                        
                                        compress_module compress_596 (
                                            .x(u[2][84]),
                                            .d(10),
                                            .result(com_out[2][84])
                                        );
                                        
                                        compress_module compress_597 (
                                            .x(u[2][85]),
                                            .d(10),
                                            .result(com_out[2][85])
                                        );
                                        
                                        compress_module compress_598 (
                                            .x(u[2][86]),
                                            .d(10),
                                            .result(com_out[2][86])
                                        );
                                        
                                        compress_module compress_599 (
                                            .x(u[2][87]),
                                            .d(10),
                                            .result(com_out[2][87])
                                        );
                                        
                                        compress_module compress_600 (
                                            .x(u[2][88]),
                                            .d(10),
                                            .result(com_out[2][88])
                                        );
                                        
                                        compress_module compress_601 (
                                            .x(u[2][89]),
                                            .d(10),
                                            .result(com_out[2][89])
                                        );
                                        
                                        compress_module compress_602 (
                                            .x(u[2][90]),
                                            .d(10),
                                            .result(com_out[2][90])
                                        );
                                        
                                        compress_module compress_603 (
                                            .x(u[2][91]),
                                            .d(10),
                                            .result(com_out[2][91])
                                        );
                                        
                                        compress_module compress_604 (
                                            .x(u[2][92]),
                                            .d(10),
                                            .result(com_out[2][92])
                                        );
                                        
                                        compress_module compress_605 (
                                            .x(u[2][93]),
                                            .d(10),
                                            .result(com_out[2][93])
                                        );
                                        
                                        compress_module compress_606 (
                                            .x(u[2][94]),
                                            .d(10),
                                            .result(com_out[2][94])
                                        );
                                        
                                        compress_module compress_607 (
                                            .x(u[2][95]),
                                            .d(10),
                                            .result(com_out[2][95])
                                        );
                                        
                                        compress_module compress_608 (
                                            .x(u[2][96]),
                                            .d(10),
                                            .result(com_out[2][96])
                                        );
                                        
                                        compress_module compress_609 (
                                            .x(u[2][97]),
                                            .d(10),
                                            .result(com_out[2][97])
                                        );
                                        
                                        compress_module compress_610 (
                                            .x(u[2][98]),
                                            .d(10),
                                            .result(com_out[2][98])
                                        );
                                        
                                        compress_module compress_611 (
                                            .x(u[2][99]),
                                            .d(10),
                                            .result(com_out[2][99])
                                        );
                                        
                                        compress_module compress_612 (
                                            .x(u[2][100]),
                                            .d(10),
                                            .result(com_out[2][100])
                                        );
                                        
                                        compress_module compress_613 (
                                            .x(u[2][101]),
                                            .d(10),
                                            .result(com_out[2][101])
                                        );
                                        
                                        compress_module compress_614 (
                                            .x(u[2][102]),
                                            .d(10),
                                            .result(com_out[2][102])
                                        );
                                        
                                        compress_module compress_615 (
                                            .x(u[2][103]),
                                            .d(10),
                                            .result(com_out[2][103])
                                        );
                                        
                                        compress_module compress_616 (
                                            .x(u[2][104]),
                                            .d(10),
                                            .result(com_out[2][104])
                                        );
                                        
                                        compress_module compress_617 (
                                            .x(u[2][105]),
                                            .d(10),
                                            .result(com_out[2][105])
                                        );
                                        
                                        compress_module compress_618 (
                                            .x(u[2][106]),
                                            .d(10),
                                            .result(com_out[2][106])
                                        );
                                        
                                        compress_module compress_619 (
                                            .x(u[2][107]),
                                            .d(10),
                                            .result(com_out[2][107])
                                        );
                                        
                                        compress_module compress_620 (
                                            .x(u[2][108]),
                                            .d(10),
                                            .result(com_out[2][108])
                                        );
                                        
                                        compress_module compress_621 (
                                            .x(u[2][109]),
                                            .d(10),
                                            .result(com_out[2][109])
                                        );
                                        
                                        compress_module compress_622 (
                                            .x(u[2][110]),
                                            .d(10),
                                            .result(com_out[2][110])
                                        );
                                        
                                        compress_module compress_623 (
                                            .x(u[2][111]),
                                            .d(10),
                                            .result(com_out[2][111])
                                        );
                                        
                                        compress_module compress_624 (
                                            .x(u[2][112]),
                                            .d(10),
                                            .result(com_out[2][112])
                                        );
                                        
                                        compress_module compress_625 (
                                            .x(u[2][113]),
                                            .d(10),
                                            .result(com_out[2][113])
                                        );
                                        
                                        compress_module compress_626 (
                                            .x(u[2][114]),
                                            .d(10),
                                            .result(com_out[2][114])
                                        );
                                        
                                        compress_module compress_627 (
                                            .x(u[2][115]),
                                            .d(10),
                                            .result(com_out[2][115])
                                        );
                                        
                                        compress_module compress_628 (
                                            .x(u[2][116]),
                                            .d(10),
                                            .result(com_out[2][116])
                                        );
                                        
                                        compress_module compress_629 (
                                            .x(u[2][117]),
                                            .d(10),
                                            .result(com_out[2][117])
                                        );
                                        
                                        compress_module compress_630 (
                                            .x(u[2][118]),
                                            .d(10),
                                            .result(com_out[2][118])
                                        );
                                        
                                        compress_module compress_631 (
                                            .x(u[2][119]),
                                            .d(10),
                                            .result(com_out[2][119])
                                        );
                                        
                                        compress_module compress_632 (
                                            .x(u[2][120]),
                                            .d(10),
                                            .result(com_out[2][120])
                                        );
                                        
                                        compress_module compress_633 (
                                            .x(u[2][121]),
                                            .d(10),
                                            .result(com_out[2][121])
                                        );
                                        
                                        compress_module compress_634 (
                                            .x(u[2][122]),
                                            .d(10),
                                            .result(com_out[2][122])
                                        );
                                        
                                        compress_module compress_635 (
                                            .x(u[2][123]),
                                            .d(10),
                                            .result(com_out[2][123])
                                        );
                                        
                                        compress_module compress_636 (
                                            .x(u[2][124]),
                                            .d(10),
                                            .result(com_out[2][124])
                                        );
                                        
                                        compress_module compress_637 (
                                            .x(u[2][125]),
                                            .d(10),
                                            .result(com_out[2][125])
                                        );
                                        
                                        compress_module compress_638 (
                                            .x(u[2][126]),
                                            .d(10),
                                            .result(com_out[2][126])
                                        );
                                        
                                        compress_module compress_639 (
                                            .x(u[2][127]),
                                            .d(10),
                                            .result(com_out[2][127])
                                        );
                                        
                                        compress_module compress_640 (
                                            .x(u[2][128]),
                                            .d(10),
                                            .result(com_out[2][128])
                                        );
                                        
                                        compress_module compress_641 (
                                            .x(u[2][129]),
                                            .d(10),
                                            .result(com_out[2][129])
                                        );
                                        
                                        compress_module compress_642 (
                                            .x(u[2][130]),
                                            .d(10),
                                            .result(com_out[2][130])
                                        );
                                        
                                        compress_module compress_643 (
                                            .x(u[2][131]),
                                            .d(10),
                                            .result(com_out[2][131])
                                        );
                                        
                                        compress_module compress_644 (
                                            .x(u[2][132]),
                                            .d(10),
                                            .result(com_out[2][132])
                                        );
                                        
                                        compress_module compress_645 (
                                            .x(u[2][133]),
                                            .d(10),
                                            .result(com_out[2][133])
                                        );
                                        
                                        compress_module compress_646 (
                                            .x(u[2][134]),
                                            .d(10),
                                            .result(com_out[2][134])
                                        );
                                        
                                        compress_module compress_647 (
                                            .x(u[2][135]),
                                            .d(10),
                                            .result(com_out[2][135])
                                        );
                                        
                                        compress_module compress_648 (
                                            .x(u[2][136]),
                                            .d(10),
                                            .result(com_out[2][136])
                                        );
                                        
                                        compress_module compress_649 (
                                            .x(u[2][137]),
                                            .d(10),
                                            .result(com_out[2][137])
                                        );
                                        
                                        compress_module compress_650 (
                                            .x(u[2][138]),
                                            .d(10),
                                            .result(com_out[2][138])
                                        );
                                        
                                        compress_module compress_651 (
                                            .x(u[2][139]),
                                            .d(10),
                                            .result(com_out[2][139])
                                        );
                                        
                                        compress_module compress_652 (
                                            .x(u[2][140]),
                                            .d(10),
                                            .result(com_out[2][140])
                                        );
                                        
                                        compress_module compress_653 (
                                            .x(u[2][141]),
                                            .d(10),
                                            .result(com_out[2][141])
                                        );
                                        
                                        compress_module compress_654 (
                                            .x(u[2][142]),
                                            .d(10),
                                            .result(com_out[2][142])
                                        );
                                        
                                        compress_module compress_655 (
                                            .x(u[2][143]),
                                            .d(10),
                                            .result(com_out[2][143])
                                        );
                                        
                                        compress_module compress_656 (
                                            .x(u[2][144]),
                                            .d(10),
                                            .result(com_out[2][144])
                                        );
                                        
                                        compress_module compress_657 (
                                            .x(u[2][145]),
                                            .d(10),
                                            .result(com_out[2][145])
                                        );
                                        
                                        compress_module compress_658 (
                                            .x(u[2][146]),
                                            .d(10),
                                            .result(com_out[2][146])
                                        );
                                        
                                        compress_module compress_659 (
                                            .x(u[2][147]),
                                            .d(10),
                                            .result(com_out[2][147])
                                        );
                                        
                                        compress_module compress_660 (
                                            .x(u[2][148]),
                                            .d(10),
                                            .result(com_out[2][148])
                                        );
                                        
                                        compress_module compress_661 (
                                            .x(u[2][149]),
                                            .d(10),
                                            .result(com_out[2][149])
                                        );
                                        
                                        compress_module compress_662 (
                                            .x(u[2][150]),
                                            .d(10),
                                            .result(com_out[2][150])
                                        );
                                        
                                        compress_module compress_663 (
                                            .x(u[2][151]),
                                            .d(10),
                                            .result(com_out[2][151])
                                        );
                                        
                                        compress_module compress_664 (
                                            .x(u[2][152]),
                                            .d(10),
                                            .result(com_out[2][152])
                                        );
                                        
                                        compress_module compress_665 (
                                            .x(u[2][153]),
                                            .d(10),
                                            .result(com_out[2][153])
                                        );
                                        
                                        compress_module compress_666 (
                                            .x(u[2][154]),
                                            .d(10),
                                            .result(com_out[2][154])
                                        );
                                        
                                        compress_module compress_667 (
                                            .x(u[2][155]),
                                            .d(10),
                                            .result(com_out[2][155])
                                        );
                                        
                                        compress_module compress_668 (
                                            .x(u[2][156]),
                                            .d(10),
                                            .result(com_out[2][156])
                                        );
                                        
                                        compress_module compress_669 (
                                            .x(u[2][157]),
                                            .d(10),
                                            .result(com_out[2][157])
                                        );
                                        
                                        compress_module compress_670 (
                                            .x(u[2][158]),
                                            .d(10),
                                            .result(com_out[2][158])
                                        );
                                        
                                        compress_module compress_671 (
                                            .x(u[2][159]),
                                            .d(10),
                                            .result(com_out[2][159])
                                        );
                                        
                                        compress_module compress_672 (
                                            .x(u[2][160]),
                                            .d(10),
                                            .result(com_out[2][160])
                                        );
                                        
                                        compress_module compress_673 (
                                            .x(u[2][161]),
                                            .d(10),
                                            .result(com_out[2][161])
                                        );
                                        
                                        compress_module compress_674 (
                                            .x(u[2][162]),
                                            .d(10),
                                            .result(com_out[2][162])
                                        );
                                        
                                        compress_module compress_675 (
                                            .x(u[2][163]),
                                            .d(10),
                                            .result(com_out[2][163])
                                        );
                                        
                                        compress_module compress_676 (
                                            .x(u[2][164]),
                                            .d(10),
                                            .result(com_out[2][164])
                                        );
                                        
                                        compress_module compress_677 (
                                            .x(u[2][165]),
                                            .d(10),
                                            .result(com_out[2][165])
                                        );
                                        
                                        compress_module compress_678 (
                                            .x(u[2][166]),
                                            .d(10),
                                            .result(com_out[2][166])
                                        );
                                        
                                        compress_module compress_679 (
                                            .x(u[2][167]),
                                            .d(10),
                                            .result(com_out[2][167])
                                        );
                                        
                                        compress_module compress_680 (
                                            .x(u[2][168]),
                                            .d(10),
                                            .result(com_out[2][168])
                                        );
                                        
                                        compress_module compress_681 (
                                            .x(u[2][169]),
                                            .d(10),
                                            .result(com_out[2][169])
                                        );
                                        
                                        compress_module compress_682 (
                                            .x(u[2][170]),
                                            .d(10),
                                            .result(com_out[2][170])
                                        );
                                        
                                        compress_module compress_683 (
                                            .x(u[2][171]),
                                            .d(10),
                                            .result(com_out[2][171])
                                        );
                                        
                                        compress_module compress_684 (
                                            .x(u[2][172]),
                                            .d(10),
                                            .result(com_out[2][172])
                                        );
                                        
                                        compress_module compress_685 (
                                            .x(u[2][173]),
                                            .d(10),
                                            .result(com_out[2][173])
                                        );
                                        
                                        compress_module compress_686 (
                                            .x(u[2][174]),
                                            .d(10),
                                            .result(com_out[2][174])
                                        );
                                        
                                        compress_module compress_687 (
                                            .x(u[2][175]),
                                            .d(10),
                                            .result(com_out[2][175])
                                        );
                                        
                                        compress_module compress_688 (
                                            .x(u[2][176]),
                                            .d(10),
                                            .result(com_out[2][176])
                                        );
                                        
                                        compress_module compress_689 (
                                            .x(u[2][177]),
                                            .d(10),
                                            .result(com_out[2][177])
                                        );
                                        
                                        compress_module compress_690 (
                                            .x(u[2][178]),
                                            .d(10),
                                            .result(com_out[2][178])
                                        );
                                        
                                        compress_module compress_691 (
                                            .x(u[2][179]),
                                            .d(10),
                                            .result(com_out[2][179])
                                        );
                                        
                                        compress_module compress_692 (
                                            .x(u[2][180]),
                                            .d(10),
                                            .result(com_out[2][180])
                                        );
                                        
                                        compress_module compress_693 (
                                            .x(u[2][181]),
                                            .d(10),
                                            .result(com_out[2][181])
                                        );
                                        
                                        compress_module compress_694 (
                                            .x(u[2][182]),
                                            .d(10),
                                            .result(com_out[2][182])
                                        );
                                        
                                        compress_module compress_695 (
                                            .x(u[2][183]),
                                            .d(10),
                                            .result(com_out[2][183])
                                        );
                                        
                                        compress_module compress_696 (
                                            .x(u[2][184]),
                                            .d(10),
                                            .result(com_out[2][184])
                                        );
                                        
                                        compress_module compress_697 (
                                            .x(u[2][185]),
                                            .d(10),
                                            .result(com_out[2][185])
                                        );
                                        
                                        compress_module compress_698 (
                                            .x(u[2][186]),
                                            .d(10),
                                            .result(com_out[2][186])
                                        );
                                        
                                        compress_module compress_699 (
                                            .x(u[2][187]),
                                            .d(10),
                                            .result(com_out[2][187])
                                        );
                                        
                                        compress_module compress_700 (
                                            .x(u[2][188]),
                                            .d(10),
                                            .result(com_out[2][188])
                                        );
                                        
                                        compress_module compress_701 (
                                            .x(u[2][189]),
                                            .d(10),
                                            .result(com_out[2][189])
                                        );
                                        
                                        compress_module compress_702 (
                                            .x(u[2][190]),
                                            .d(10),
                                            .result(com_out[2][190])
                                        );
                                        
                                        compress_module compress_703 (
                                            .x(u[2][191]),
                                            .d(10),
                                            .result(com_out[2][191])
                                        );
                                        
                                        compress_module compress_704 (
                                            .x(u[2][192]),
                                            .d(10),
                                            .result(com_out[2][192])
                                        );
                                        
                                        compress_module compress_705 (
                                            .x(u[2][193]),
                                            .d(10),
                                            .result(com_out[2][193])
                                        );
                                        
                                        compress_module compress_706 (
                                            .x(u[2][194]),
                                            .d(10),
                                            .result(com_out[2][194])
                                        );
                                        
                                        compress_module compress_707 (
                                            .x(u[2][195]),
                                            .d(10),
                                            .result(com_out[2][195])
                                        );
                                        
                                        compress_module compress_708 (
                                            .x(u[2][196]),
                                            .d(10),
                                            .result(com_out[2][196])
                                        );
                                        
                                        compress_module compress_709 (
                                            .x(u[2][197]),
                                            .d(10),
                                            .result(com_out[2][197])
                                        );
                                        
                                        compress_module compress_710 (
                                            .x(u[2][198]),
                                            .d(10),
                                            .result(com_out[2][198])
                                        );
                                        
                                        compress_module compress_711 (
                                            .x(u[2][199]),
                                            .d(10),
                                            .result(com_out[2][199])
                                        );
                                        
                                        compress_module compress_712 (
                                            .x(u[2][200]),
                                            .d(10),
                                            .result(com_out[2][200])
                                        );
                                        
                                        compress_module compress_713 (
                                            .x(u[2][201]),
                                            .d(10),
                                            .result(com_out[2][201])
                                        );
                                        
                                        compress_module compress_714 (
                                            .x(u[2][202]),
                                            .d(10),
                                            .result(com_out[2][202])
                                        );
                                        
                                        compress_module compress_715 (
                                            .x(u[2][203]),
                                            .d(10),
                                            .result(com_out[2][203])
                                        );
                                        
                                        compress_module compress_716 (
                                            .x(u[2][204]),
                                            .d(10),
                                            .result(com_out[2][204])
                                        );
                                        
                                        compress_module compress_717 (
                                            .x(u[2][205]),
                                            .d(10),
                                            .result(com_out[2][205])
                                        );
                                        
                                        compress_module compress_718 (
                                            .x(u[2][206]),
                                            .d(10),
                                            .result(com_out[2][206])
                                        );
                                        
                                        compress_module compress_719 (
                                            .x(u[2][207]),
                                            .d(10),
                                            .result(com_out[2][207])
                                        );
                                        
                                        compress_module compress_720 (
                                            .x(u[2][208]),
                                            .d(10),
                                            .result(com_out[2][208])
                                        );
                                        
                                        compress_module compress_721 (
                                            .x(u[2][209]),
                                            .d(10),
                                            .result(com_out[2][209])
                                        );
                                        
                                        compress_module compress_722 (
                                            .x(u[2][210]),
                                            .d(10),
                                            .result(com_out[2][210])
                                        );
                                        
                                        compress_module compress_723 (
                                            .x(u[2][211]),
                                            .d(10),
                                            .result(com_out[2][211])
                                        );
                                        
                                        compress_module compress_724 (
                                            .x(u[2][212]),
                                            .d(10),
                                            .result(com_out[2][212])
                                        );
                                        
                                        compress_module compress_725 (
                                            .x(u[2][213]),
                                            .d(10),
                                            .result(com_out[2][213])
                                        );
                                        
                                        compress_module compress_726 (
                                            .x(u[2][214]),
                                            .d(10),
                                            .result(com_out[2][214])
                                        );
                                        
                                        compress_module compress_727 (
                                            .x(u[2][215]),
                                            .d(10),
                                            .result(com_out[2][215])
                                        );
                                        
                                        compress_module compress_728 (
                                            .x(u[2][216]),
                                            .d(10),
                                            .result(com_out[2][216])
                                        );
                                        
                                        compress_module compress_729 (
                                            .x(u[2][217]),
                                            .d(10),
                                            .result(com_out[2][217])
                                        );
                                        
                                        compress_module compress_730 (
                                            .x(u[2][218]),
                                            .d(10),
                                            .result(com_out[2][218])
                                        );
                                        
                                        compress_module compress_731 (
                                            .x(u[2][219]),
                                            .d(10),
                                            .result(com_out[2][219])
                                        );
                                        
                                        compress_module compress_732 (
                                            .x(u[2][220]),
                                            .d(10),
                                            .result(com_out[2][220])
                                        );
                                        
                                        compress_module compress_733 (
                                            .x(u[2][221]),
                                            .d(10),
                                            .result(com_out[2][221])
                                        );
                                        
                                        compress_module compress_734 (
                                            .x(u[2][222]),
                                            .d(10),
                                            .result(com_out[2][222])
                                        );
                                        
                                        compress_module compress_735 (
                                            .x(u[2][223]),
                                            .d(10),
                                            .result(com_out[2][223])
                                        );
                                        
                                        compress_module compress_736 (
                                            .x(u[2][224]),
                                            .d(10),
                                            .result(com_out[2][224])
                                        );
                                        
                                        compress_module compress_737 (
                                            .x(u[2][225]),
                                            .d(10),
                                            .result(com_out[2][225])
                                        );
                                        
                                        compress_module compress_738 (
                                            .x(u[2][226]),
                                            .d(10),
                                            .result(com_out[2][226])
                                        );
                                        
                                        compress_module compress_739 (
                                            .x(u[2][227]),
                                            .d(10),
                                            .result(com_out[2][227])
                                        );
                                        
                                        compress_module compress_740 (
                                            .x(u[2][228]),
                                            .d(10),
                                            .result(com_out[2][228])
                                        );
                                        
                                        compress_module compress_741 (
                                            .x(u[2][229]),
                                            .d(10),
                                            .result(com_out[2][229])
                                        );
                                        
                                        compress_module compress_742 (
                                            .x(u[2][230]),
                                            .d(10),
                                            .result(com_out[2][230])
                                        );
                                        
                                        compress_module compress_743 (
                                            .x(u[2][231]),
                                            .d(10),
                                            .result(com_out[2][231])
                                        );
                                        
                                        compress_module compress_744 (
                                            .x(u[2][232]),
                                            .d(10),
                                            .result(com_out[2][232])
                                        );
                                        
                                        compress_module compress_745 (
                                            .x(u[2][233]),
                                            .d(10),
                                            .result(com_out[2][233])
                                        );
                                        
                                        compress_module compress_746 (
                                            .x(u[2][234]),
                                            .d(10),
                                            .result(com_out[2][234])
                                        );
                                        
                                        compress_module compress_747 (
                                            .x(u[2][235]),
                                            .d(10),
                                            .result(com_out[2][235])
                                        );
                                        
                                        compress_module compress_748 (
                                            .x(u[2][236]),
                                            .d(10),
                                            .result(com_out[2][236])
                                        );
                                        
                                        compress_module compress_749 (
                                            .x(u[2][237]),
                                            .d(10),
                                            .result(com_out[2][237])
                                        );
                                        
                                        compress_module compress_750 (
                                            .x(u[2][238]),
                                            .d(10),
                                            .result(com_out[2][238])
                                        );
                                        
                                        compress_module compress_751 (
                                            .x(u[2][239]),
                                            .d(10),
                                            .result(com_out[2][239])
                                        );
                                        
                                        compress_module compress_752 (
                                            .x(u[2][240]),
                                            .d(10),
                                            .result(com_out[2][240])
                                        );
                                        
                                        compress_module compress_753 (
                                            .x(u[2][241]),
                                            .d(10),
                                            .result(com_out[2][241])
                                        );
                                        
                                        compress_module compress_754 (
                                            .x(u[2][242]),
                                            .d(10),
                                            .result(com_out[2][242])
                                        );
                                        
                                        compress_module compress_755 (
                                            .x(u[2][243]),
                                            .d(10),
                                            .result(com_out[2][243])
                                        );
                                        
                                        compress_module compress_756 (
                                            .x(u[2][244]),
                                            .d(10),
                                            .result(com_out[2][244])
                                        );
                                        
                                        compress_module compress_757 (
                                            .x(u[2][245]),
                                            .d(10),
                                            .result(com_out[2][245])
                                        );
                                        
                                        compress_module compress_758 (
                                            .x(u[2][246]),
                                            .d(10),
                                            .result(com_out[2][246])
                                        );
                                        
                                        compress_module compress_759 (
                                            .x(u[2][247]),
                                            .d(10),
                                            .result(com_out[2][247])
                                        );
                                        
                                        compress_module compress_760 (
                                            .x(u[2][248]),
                                            .d(10),
                                            .result(com_out[2][248])
                                        );
                                        
                                        compress_module compress_761 (
                                            .x(u[2][249]),
                                            .d(10),
                                            .result(com_out[2][249])
                                        );
                                        
                                        compress_module compress_762 (
                                            .x(u[2][250]),
                                            .d(10),
                                            .result(com_out[2][250])
                                        );
                                        
                                        compress_module compress_763 (
                                            .x(u[2][251]),
                                            .d(10),
                                            .result(com_out[2][251])
                                        );
                                        
                                        compress_module compress_764 (
                                            .x(u[2][252]),
                                            .d(10),
                                            .result(com_out[2][252])
                                        );
                                        
                                        compress_module compress_765 (
                                            .x(u[2][253]),
                                            .d(10),
                                            .result(com_out[2][253])
                                        );
                                        
                                        compress_module compress_766 (
                                            .x(u[2][254]),
                                            .d(10),
                                            .result(com_out[2][254])
                                        );
                                        
                                        compress_module compress_767 (
                                            .x(u[2][255]),
                                            .d(10),
                                            .result(com_out[2][255])
                                        );
                                        compress_module comp_v_0 (
                                            .x(result[0][0]),
                                            .d(4),
                                            .result(comp_v[0][0])
                                        );
                                        
                                        compress_module comp_v_1 (
                                            .x(result[0][1]),
                                            .d(4),
                                            .result(comp_v[0][1])
                                        );
                                        
                                        compress_module comp_v_2 (
                                            .x(result[0][2]),
                                            .d(4),
                                            .result(comp_v[0][2])
                                        );
                                        
                                        compress_module comp_v_3 (
                                            .x(result[0][3]),
                                            .d(4),
                                            .result(comp_v[0][3])
                                        );
                                        
                                        compress_module comp_v_4 (
                                            .x(result[0][4]),
                                            .d(4),
                                            .result(comp_v[0][4])
                                        );
                                        
                                        compress_module comp_v_5 (
                                            .x(result[0][5]),
                                            .d(4),
                                            .result(comp_v[0][5])
                                        );
                                        
                                        compress_module comp_v_6 (
                                            .x(result[0][6]),
                                            .d(4),
                                            .result(comp_v[0][6])
                                        );
                                        
                                        compress_module comp_v_7 (
                                            .x(result[0][7]),
                                            .d(4),
                                            .result(comp_v[0][7])
                                        );
                                        
                                        compress_module comp_v_8 (
                                            .x(result[0][8]),
                                            .d(4),
                                            .result(comp_v[0][8])
                                        );
                                        
                                        compress_module comp_v_9 (
                                            .x(result[0][9]),
                                            .d(4),
                                            .result(comp_v[0][9])
                                        );
                                        
                                        compress_module comp_v_10 (
                                            .x(result[0][10]),
                                            .d(4),
                                            .result(comp_v[0][10])
                                        );
                                        
                                        compress_module comp_v_11 (
                                            .x(result[0][11]),
                                            .d(4),
                                            .result(comp_v[0][11])
                                        );
                                        
                                        compress_module comp_v_12 (
                                            .x(result[0][12]),
                                            .d(4),
                                            .result(comp_v[0][12])
                                        );
                                        
                                        compress_module comp_v_13 (
                                            .x(result[0][13]),
                                            .d(4),
                                            .result(comp_v[0][13])
                                        );
                                        
                                        compress_module comp_v_14 (
                                            .x(result[0][14]),
                                            .d(4),
                                            .result(comp_v[0][14])
                                        );
                                        
                                        compress_module comp_v_15 (
                                            .x(result[0][15]),
                                            .d(4),
                                            .result(comp_v[0][15])
                                        );
                                        
                                        compress_module comp_v_16 (
                                            .x(result[0][16]),
                                            .d(4),
                                            .result(comp_v[0][16])
                                        );
                                        
                                        compress_module comp_v_17 (
                                            .x(result[0][17]),
                                            .d(4),
                                            .result(comp_v[0][17])
                                        );
                                        
                                        compress_module comp_v_18 (
                                            .x(result[0][18]),
                                            .d(4),
                                            .result(comp_v[0][18])
                                        );
                                        
                                        compress_module comp_v_19 (
                                            .x(result[0][19]),
                                            .d(4),
                                            .result(comp_v[0][19])
                                        );
                                        
                                        compress_module comp_v_20 (
                                            .x(result[0][20]),
                                            .d(4),
                                            .result(comp_v[0][20])
                                        );
                                        
                                        compress_module comp_v_21 (
                                            .x(result[0][21]),
                                            .d(4),
                                            .result(comp_v[0][21])
                                        );
                                        
                                        compress_module comp_v_22 (
                                            .x(result[0][22]),
                                            .d(4),
                                            .result(comp_v[0][22])
                                        );
                                        
                                        compress_module comp_v_23 (
                                            .x(result[0][23]),
                                            .d(4),
                                            .result(comp_v[0][23])
                                        );
                                        
                                        compress_module comp_v_24 (
                                            .x(result[0][24]),
                                            .d(4),
                                            .result(comp_v[0][24])
                                        );
                                        
                                        compress_module comp_v_25 (
                                            .x(result[0][25]),
                                            .d(4),
                                            .result(comp_v[0][25])
                                        );
                                        
                                        compress_module comp_v_26 (
                                            .x(result[0][26]),
                                            .d(4),
                                            .result(comp_v[0][26])
                                        );
                                        
                                        compress_module comp_v_27 (
                                            .x(result[0][27]),
                                            .d(4),
                                            .result(comp_v[0][27])
                                        );
                                        
                                        compress_module comp_v_28 (
                                            .x(result[0][28]),
                                            .d(4),
                                            .result(comp_v[0][28])
                                        );
                                        
                                        compress_module comp_v_29 (
                                            .x(result[0][29]),
                                            .d(4),
                                            .result(comp_v[0][29])
                                        );
                                        
                                        compress_module comp_v_30 (
                                            .x(result[0][30]),
                                            .d(4),
                                            .result(comp_v[0][30])
                                        );
                                        
                                        compress_module comp_v_31 (
                                            .x(result[0][31]),
                                            .d(4),
                                            .result(comp_v[0][31])
                                        );
                                        
                                        compress_module comp_v_32 (
                                            .x(result[0][32]),
                                            .d(4),
                                            .result(comp_v[0][32])
                                        );
                                        
                                        compress_module comp_v_33 (
                                            .x(result[0][33]),
                                            .d(4),
                                            .result(comp_v[0][33])
                                        );
                                        
                                        compress_module comp_v_34 (
                                            .x(result[0][34]),
                                            .d(4),
                                            .result(comp_v[0][34])
                                        );
                                        
                                        compress_module comp_v_35 (
                                            .x(result[0][35]),
                                            .d(4),
                                            .result(comp_v[0][35])
                                        );
                                        
                                        compress_module comp_v_36 (
                                            .x(result[0][36]),
                                            .d(4),
                                            .result(comp_v[0][36])
                                        );
                                        
                                        compress_module comp_v_37 (
                                            .x(result[0][37]),
                                            .d(4),
                                            .result(comp_v[0][37])
                                        );
                                        
                                        compress_module comp_v_38 (
                                            .x(result[0][38]),
                                            .d(4),
                                            .result(comp_v[0][38])
                                        );
                                        
                                        compress_module comp_v_39 (
                                            .x(result[0][39]),
                                            .d(4),
                                            .result(comp_v[0][39])
                                        );
                                        
                                        compress_module comp_v_40 (
                                            .x(result[0][40]),
                                            .d(4),
                                            .result(comp_v[0][40])
                                        );
                                        
                                        compress_module comp_v_41 (
                                            .x(result[0][41]),
                                            .d(4),
                                            .result(comp_v[0][41])
                                        );
                                        
                                        compress_module comp_v_42 (
                                            .x(result[0][42]),
                                            .d(4),
                                            .result(comp_v[0][42])
                                        );
                                        
                                        compress_module comp_v_43 (
                                            .x(result[0][43]),
                                            .d(4),
                                            .result(comp_v[0][43])
                                        );
                                        
                                        compress_module comp_v_44 (
                                            .x(result[0][44]),
                                            .d(4),
                                            .result(comp_v[0][44])
                                        );
                                        
                                        compress_module comp_v_45 (
                                            .x(result[0][45]),
                                            .d(4),
                                            .result(comp_v[0][45])
                                        );
                                        
                                        compress_module comp_v_46 (
                                            .x(result[0][46]),
                                            .d(4),
                                            .result(comp_v[0][46])
                                        );
                                        
                                        compress_module comp_v_47 (
                                            .x(result[0][47]),
                                            .d(4),
                                            .result(comp_v[0][47])
                                        );
                                        
                                        compress_module comp_v_48 (
                                            .x(result[0][48]),
                                            .d(4),
                                            .result(comp_v[0][48])
                                        );
                                        
                                        compress_module comp_v_49 (
                                            .x(result[0][49]),
                                            .d(4),
                                            .result(comp_v[0][49])
                                        );
                                        
                                        compress_module comp_v_50 (
                                            .x(result[0][50]),
                                            .d(4),
                                            .result(comp_v[0][50])
                                        );
                                        
                                        compress_module comp_v_51 (
                                            .x(result[0][51]),
                                            .d(4),
                                            .result(comp_v[0][51])
                                        );
                                        
                                        compress_module comp_v_52 (
                                            .x(result[0][52]),
                                            .d(4),
                                            .result(comp_v[0][52])
                                        );
                                        
                                        compress_module comp_v_53 (
                                            .x(result[0][53]),
                                            .d(4),
                                            .result(comp_v[0][53])
                                        );
                                        
                                        compress_module comp_v_54 (
                                            .x(result[0][54]),
                                            .d(4),
                                            .result(comp_v[0][54])
                                        );
                                        
                                        compress_module comp_v_55 (
                                            .x(result[0][55]),
                                            .d(4),
                                            .result(comp_v[0][55])
                                        );
                                        
                                        compress_module comp_v_56 (
                                            .x(result[0][56]),
                                            .d(4),
                                            .result(comp_v[0][56])
                                        );
                                        
                                        compress_module comp_v_57 (
                                            .x(result[0][57]),
                                            .d(4),
                                            .result(comp_v[0][57])
                                        );
                                        
                                        compress_module comp_v_58 (
                                            .x(result[0][58]),
                                            .d(4),
                                            .result(comp_v[0][58])
                                        );
                                        
                                        compress_module comp_v_59 (
                                            .x(result[0][59]),
                                            .d(4),
                                            .result(comp_v[0][59])
                                        );
                                        
                                        compress_module comp_v_60 (
                                            .x(result[0][60]),
                                            .d(4),
                                            .result(comp_v[0][60])
                                        );
                                        
                                        compress_module comp_v_61 (
                                            .x(result[0][61]),
                                            .d(4),
                                            .result(comp_v[0][61])
                                        );
                                        
                                        compress_module comp_v_62 (
                                            .x(result[0][62]),
                                            .d(4),
                                            .result(comp_v[0][62])
                                        );
                                        
                                        compress_module comp_v_63 (
                                            .x(result[0][63]),
                                            .d(4),
                                            .result(comp_v[0][63])
                                        );
                                        
                                        compress_module comp_v_64 (
                                            .x(result[0][64]),
                                            .d(4),
                                            .result(comp_v[0][64])
                                        );
                                        
                                        compress_module comp_v_65 (
                                            .x(result[0][65]),
                                            .d(4),
                                            .result(comp_v[0][65])
                                        );
                                        
                                        compress_module comp_v_66 (
                                            .x(result[0][66]),
                                            .d(4),
                                            .result(comp_v[0][66])
                                        );
                                        
                                        compress_module comp_v_67 (
                                            .x(result[0][67]),
                                            .d(4),
                                            .result(comp_v[0][67])
                                        );
                                        
                                        compress_module comp_v_68 (
                                            .x(result[0][68]),
                                            .d(4),
                                            .result(comp_v[0][68])
                                        );
                                        
                                        compress_module comp_v_69 (
                                            .x(result[0][69]),
                                            .d(4),
                                            .result(comp_v[0][69])
                                        );
                                        
                                        compress_module comp_v_70 (
                                            .x(result[0][70]),
                                            .d(4),
                                            .result(comp_v[0][70])
                                        );
                                        
                                        compress_module comp_v_71 (
                                            .x(result[0][71]),
                                            .d(4),
                                            .result(comp_v[0][71])
                                        );
                                        
                                        compress_module comp_v_72 (
                                            .x(result[0][72]),
                                            .d(4),
                                            .result(comp_v[0][72])
                                        );
                                        
                                        compress_module comp_v_73 (
                                            .x(result[0][73]),
                                            .d(4),
                                            .result(comp_v[0][73])
                                        );
                                        
                                        compress_module comp_v_74 (
                                            .x(result[0][74]),
                                            .d(4),
                                            .result(comp_v[0][74])
                                        );
                                        
                                        compress_module comp_v_75 (
                                            .x(result[0][75]),
                                            .d(4),
                                            .result(comp_v[0][75])
                                        );
                                        
                                        compress_module comp_v_76 (
                                            .x(result[0][76]),
                                            .d(4),
                                            .result(comp_v[0][76])
                                        );
                                        
                                        compress_module comp_v_77 (
                                            .x(result[0][77]),
                                            .d(4),
                                            .result(comp_v[0][77])
                                        );
                                        
                                        compress_module comp_v_78 (
                                            .x(result[0][78]),
                                            .d(4),
                                            .result(comp_v[0][78])
                                        );
                                        
                                        compress_module comp_v_79 (
                                            .x(result[0][79]),
                                            .d(4),
                                            .result(comp_v[0][79])
                                        );
                                        
                                        compress_module comp_v_80 (
                                            .x(result[0][80]),
                                            .d(4),
                                            .result(comp_v[0][80])
                                        );
                                        
                                        compress_module comp_v_81 (
                                            .x(result[0][81]),
                                            .d(4),
                                            .result(comp_v[0][81])
                                        );
                                        
                                        compress_module comp_v_82 (
                                            .x(result[0][82]),
                                            .d(4),
                                            .result(comp_v[0][82])
                                        );
                                        
                                        compress_module comp_v_83 (
                                            .x(result[0][83]),
                                            .d(4),
                                            .result(comp_v[0][83])
                                        );
                                        
                                        compress_module comp_v_84 (
                                            .x(result[0][84]),
                                            .d(4),
                                            .result(comp_v[0][84])
                                        );
                                        
                                        compress_module comp_v_85 (
                                            .x(result[0][85]),
                                            .d(4),
                                            .result(comp_v[0][85])
                                        );
                                        
                                        compress_module comp_v_86 (
                                            .x(result[0][86]),
                                            .d(4),
                                            .result(comp_v[0][86])
                                        );
                                        
                                        compress_module comp_v_87 (
                                            .x(result[0][87]),
                                            .d(4),
                                            .result(comp_v[0][87])
                                        );
                                        
                                        compress_module comp_v_88 (
                                            .x(result[0][88]),
                                            .d(4),
                                            .result(comp_v[0][88])
                                        );
                                        
                                        compress_module comp_v_89 (
                                            .x(result[0][89]),
                                            .d(4),
                                            .result(comp_v[0][89])
                                        );
                                        
                                        compress_module comp_v_90 (
                                            .x(result[0][90]),
                                            .d(4),
                                            .result(comp_v[0][90])
                                        );
                                        
                                        compress_module comp_v_91 (
                                            .x(result[0][91]),
                                            .d(4),
                                            .result(comp_v[0][91])
                                        );
                                        
                                        compress_module comp_v_92 (
                                            .x(result[0][92]),
                                            .d(4),
                                            .result(comp_v[0][92])
                                        );
                                        
                                        compress_module comp_v_93 (
                                            .x(result[0][93]),
                                            .d(4),
                                            .result(comp_v[0][93])
                                        );
                                        
                                        compress_module comp_v_94 (
                                            .x(result[0][94]),
                                            .d(4),
                                            .result(comp_v[0][94])
                                        );
                                        
                                        compress_module comp_v_95 (
                                            .x(result[0][95]),
                                            .d(4),
                                            .result(comp_v[0][95])
                                        );
                                        
                                        compress_module comp_v_96 (
                                            .x(result[0][96]),
                                            .d(4),
                                            .result(comp_v[0][96])
                                        );
                                        
                                        compress_module comp_v_97 (
                                            .x(result[0][97]),
                                            .d(4),
                                            .result(comp_v[0][97])
                                        );
                                        
                                        compress_module comp_v_98 (
                                            .x(result[0][98]),
                                            .d(4),
                                            .result(comp_v[0][98])
                                        );
                                        
                                        compress_module comp_v_99 (
                                            .x(result[0][99]),
                                            .d(4),
                                            .result(comp_v[0][99])
                                        );
                                        
                                        compress_module comp_v_100 (
                                            .x(result[0][100]),
                                            .d(4),
                                            .result(comp_v[0][100])
                                        );
                                        
                                        compress_module comp_v_101 (
                                            .x(result[0][101]),
                                            .d(4),
                                            .result(comp_v[0][101])
                                        );
                                        
                                        compress_module comp_v_102 (
                                            .x(result[0][102]),
                                            .d(4),
                                            .result(comp_v[0][102])
                                        );
                                        
                                        compress_module comp_v_103 (
                                            .x(result[0][103]),
                                            .d(4),
                                            .result(comp_v[0][103])
                                        );
                                        
                                        compress_module comp_v_104 (
                                            .x(result[0][104]),
                                            .d(4),
                                            .result(comp_v[0][104])
                                        );
                                        
                                        compress_module comp_v_105 (
                                            .x(result[0][105]),
                                            .d(4),
                                            .result(comp_v[0][105])
                                        );
                                        
                                        compress_module comp_v_106 (
                                            .x(result[0][106]),
                                            .d(4),
                                            .result(comp_v[0][106])
                                        );
                                        
                                        compress_module comp_v_107 (
                                            .x(result[0][107]),
                                            .d(4),
                                            .result(comp_v[0][107])
                                        );
                                        
                                        compress_module comp_v_108 (
                                            .x(result[0][108]),
                                            .d(4),
                                            .result(comp_v[0][108])
                                        );
                                        
                                        compress_module comp_v_109 (
                                            .x(result[0][109]),
                                            .d(4),
                                            .result(comp_v[0][109])
                                        );
                                        
                                        compress_module comp_v_110 (
                                            .x(result[0][110]),
                                            .d(4),
                                            .result(comp_v[0][110])
                                        );
                                        
                                        compress_module comp_v_111 (
                                            .x(result[0][111]),
                                            .d(4),
                                            .result(comp_v[0][111])
                                        );
                                        
                                        compress_module comp_v_112 (
                                            .x(result[0][112]),
                                            .d(4),
                                            .result(comp_v[0][112])
                                        );
                                        
                                        compress_module comp_v_113 (
                                            .x(result[0][113]),
                                            .d(4),
                                            .result(comp_v[0][113])
                                        );
                                        
                                        compress_module comp_v_114 (
                                            .x(result[0][114]),
                                            .d(4),
                                            .result(comp_v[0][114])
                                        );
                                        
                                        compress_module comp_v_115 (
                                            .x(result[0][115]),
                                            .d(4),
                                            .result(comp_v[0][115])
                                        );
                                        
                                        compress_module comp_v_116 (
                                            .x(result[0][116]),
                                            .d(4),
                                            .result(comp_v[0][116])
                                        );
                                        
                                        compress_module comp_v_117 (
                                            .x(result[0][117]),
                                            .d(4),
                                            .result(comp_v[0][117])
                                        );
                                        
                                        compress_module comp_v_118 (
                                            .x(result[0][118]),
                                            .d(4),
                                            .result(comp_v[0][118])
                                        );
                                        
                                        compress_module comp_v_119 (
                                            .x(result[0][119]),
                                            .d(4),
                                            .result(comp_v[0][119])
                                        );
                                        
                                        compress_module comp_v_120 (
                                            .x(result[0][120]),
                                            .d(4),
                                            .result(comp_v[0][120])
                                        );
                                        
                                        compress_module comp_v_121 (
                                            .x(result[0][121]),
                                            .d(4),
                                            .result(comp_v[0][121])
                                        );
                                        
                                        compress_module comp_v_122 (
                                            .x(result[0][122]),
                                            .d(4),
                                            .result(comp_v[0][122])
                                        );
                                        
                                        compress_module comp_v_123 (
                                            .x(result[0][123]),
                                            .d(4),
                                            .result(comp_v[0][123])
                                        );
                                        
                                        compress_module comp_v_124 (
                                            .x(result[0][124]),
                                            .d(4),
                                            .result(comp_v[0][124])
                                        );
                                        
                                        compress_module comp_v_125 (
                                            .x(result[0][125]),
                                            .d(4),
                                            .result(comp_v[0][125])
                                        );
                                        
                                        compress_module comp_v_126 (
                                            .x(result[0][126]),
                                            .d(4),
                                            .result(comp_v[0][126])
                                        );
                                        
                                        compress_module comp_v_127 (
                                            .x(result[0][127]),
                                            .d(4),
                                            .result(comp_v[0][127])
                                        );
                                        
                                        compress_module comp_v_128 (
                                            .x(result[0][128]),
                                            .d(4),
                                            .result(comp_v[0][128])
                                        );
                                        
                                        compress_module comp_v_129 (
                                            .x(result[0][129]),
                                            .d(4),
                                            .result(comp_v[0][129])
                                        );
                                        
                                        compress_module comp_v_130 (
                                            .x(result[0][130]),
                                            .d(4),
                                            .result(comp_v[0][130])
                                        );
                                        
                                        compress_module comp_v_131 (
                                            .x(result[0][131]),
                                            .d(4),
                                            .result(comp_v[0][131])
                                        );
                                        
                                        compress_module comp_v_132 (
                                            .x(result[0][132]),
                                            .d(4),
                                            .result(comp_v[0][132])
                                        );
                                        
                                        compress_module comp_v_133 (
                                            .x(result[0][133]),
                                            .d(4),
                                            .result(comp_v[0][133])
                                        );
                                        
                                        compress_module comp_v_134 (
                                            .x(result[0][134]),
                                            .d(4),
                                            .result(comp_v[0][134])
                                        );
                                        
                                        compress_module comp_v_135 (
                                            .x(result[0][135]),
                                            .d(4),
                                            .result(comp_v[0][135])
                                        );
                                        
                                        compress_module comp_v_136 (
                                            .x(result[0][136]),
                                            .d(4),
                                            .result(comp_v[0][136])
                                        );
                                        
                                        compress_module comp_v_137 (
                                            .x(result[0][137]),
                                            .d(4),
                                            .result(comp_v[0][137])
                                        );
                                        
                                        compress_module comp_v_138 (
                                            .x(result[0][138]),
                                            .d(4),
                                            .result(comp_v[0][138])
                                        );
                                        
                                        compress_module comp_v_139 (
                                            .x(result[0][139]),
                                            .d(4),
                                            .result(comp_v[0][139])
                                        );
                                        
                                        compress_module comp_v_140 (
                                            .x(result[0][140]),
                                            .d(4),
                                            .result(comp_v[0][140])
                                        );
                                        
                                        compress_module comp_v_141 (
                                            .x(result[0][141]),
                                            .d(4),
                                            .result(comp_v[0][141])
                                        );
                                        
                                        compress_module comp_v_142 (
                                            .x(result[0][142]),
                                            .d(4),
                                            .result(comp_v[0][142])
                                        );
                                        
                                        compress_module comp_v_143 (
                                            .x(result[0][143]),
                                            .d(4),
                                            .result(comp_v[0][143])
                                        );
                                        
                                        compress_module comp_v_144 (
                                            .x(result[0][144]),
                                            .d(4),
                                            .result(comp_v[0][144])
                                        );
                                        
                                        compress_module comp_v_145 (
                                            .x(result[0][145]),
                                            .d(4),
                                            .result(comp_v[0][145])
                                        );
                                        
                                        compress_module comp_v_146 (
                                            .x(result[0][146]),
                                            .d(4),
                                            .result(comp_v[0][146])
                                        );
                                        
                                        compress_module comp_v_147 (
                                            .x(result[0][147]),
                                            .d(4),
                                            .result(comp_v[0][147])
                                        );
                                        
                                        compress_module comp_v_148 (
                                            .x(result[0][148]),
                                            .d(4),
                                            .result(comp_v[0][148])
                                        );
                                        
                                        compress_module comp_v_149 (
                                            .x(result[0][149]),
                                            .d(4),
                                            .result(comp_v[0][149])
                                        );
                                        
                                        compress_module comp_v_150 (
                                            .x(result[0][150]),
                                            .d(4),
                                            .result(comp_v[0][150])
                                        );
                                        
                                        compress_module comp_v_151 (
                                            .x(result[0][151]),
                                            .d(4),
                                            .result(comp_v[0][151])
                                        );
                                        
                                        compress_module comp_v_152 (
                                            .x(result[0][152]),
                                            .d(4),
                                            .result(comp_v[0][152])
                                        );
                                        
                                        compress_module comp_v_153 (
                                            .x(result[0][153]),
                                            .d(4),
                                            .result(comp_v[0][153])
                                        );
                                        
                                        compress_module comp_v_154 (
                                            .x(result[0][154]),
                                            .d(4),
                                            .result(comp_v[0][154])
                                        );
                                        
                                        compress_module comp_v_155 (
                                            .x(result[0][155]),
                                            .d(4),
                                            .result(comp_v[0][155])
                                        );
                                        
                                        compress_module comp_v_156 (
                                            .x(result[0][156]),
                                            .d(4),
                                            .result(comp_v[0][156])
                                        );
                                        
                                        compress_module comp_v_157 (
                                            .x(result[0][157]),
                                            .d(4),
                                            .result(comp_v[0][157])
                                        );
                                        
                                        compress_module comp_v_158 (
                                            .x(result[0][158]),
                                            .d(4),
                                            .result(comp_v[0][158])
                                        );
                                        
                                        compress_module comp_v_159 (
                                            .x(result[0][159]),
                                            .d(4),
                                            .result(comp_v[0][159])
                                        );
                                        
                                        compress_module comp_v_160 (
                                            .x(result[0][160]),
                                            .d(4),
                                            .result(comp_v[0][160])
                                        );
                                        
                                        compress_module comp_v_161 (
                                            .x(result[0][161]),
                                            .d(4),
                                            .result(comp_v[0][161])
                                        );
                                        
                                        compress_module comp_v_162 (
                                            .x(result[0][162]),
                                            .d(4),
                                            .result(comp_v[0][162])
                                        );
                                        
                                        compress_module comp_v_163 (
                                            .x(result[0][163]),
                                            .d(4),
                                            .result(comp_v[0][163])
                                        );
                                        
                                        compress_module comp_v_164 (
                                            .x(result[0][164]),
                                            .d(4),
                                            .result(comp_v[0][164])
                                        );
                                        
                                        compress_module comp_v_165 (
                                            .x(result[0][165]),
                                            .d(4),
                                            .result(comp_v[0][165])
                                        );
                                        
                                        compress_module comp_v_166 (
                                            .x(result[0][166]),
                                            .d(4),
                                            .result(comp_v[0][166])
                                        );
                                        
                                        compress_module comp_v_167 (
                                            .x(result[0][167]),
                                            .d(4),
                                            .result(comp_v[0][167])
                                        );
                                        
                                        compress_module comp_v_168 (
                                            .x(result[0][168]),
                                            .d(4),
                                            .result(comp_v[0][168])
                                        );
                                        
                                        compress_module comp_v_169 (
                                            .x(result[0][169]),
                                            .d(4),
                                            .result(comp_v[0][169])
                                        );
                                        
                                        compress_module comp_v_170 (
                                            .x(result[0][170]),
                                            .d(4),
                                            .result(comp_v[0][170])
                                        );
                                        
                                        compress_module comp_v_171 (
                                            .x(result[0][171]),
                                            .d(4),
                                            .result(comp_v[0][171])
                                        );
                                        
                                        compress_module comp_v_172 (
                                            .x(result[0][172]),
                                            .d(4),
                                            .result(comp_v[0][172])
                                        );
                                        
                                        compress_module comp_v_173 (
                                            .x(result[0][173]),
                                            .d(4),
                                            .result(comp_v[0][173])
                                        );
                                        
                                        compress_module comp_v_174 (
                                            .x(result[0][174]),
                                            .d(4),
                                            .result(comp_v[0][174])
                                        );
                                        
                                        compress_module comp_v_175 (
                                            .x(result[0][175]),
                                            .d(4),
                                            .result(comp_v[0][175])
                                        );
                                        
                                        compress_module comp_v_176 (
                                            .x(result[0][176]),
                                            .d(4),
                                            .result(comp_v[0][176])
                                        );
                                        
                                        compress_module comp_v_177 (
                                            .x(result[0][177]),
                                            .d(4),
                                            .result(comp_v[0][177])
                                        );
                                        
                                        compress_module comp_v_178 (
                                            .x(result[0][178]),
                                            .d(4),
                                            .result(comp_v[0][178])
                                        );
                                        
                                        compress_module comp_v_179 (
                                            .x(result[0][179]),
                                            .d(4),
                                            .result(comp_v[0][179])
                                        );
                                        
                                        compress_module comp_v_180 (
                                            .x(result[0][180]),
                                            .d(4),
                                            .result(comp_v[0][180])
                                        );
                                        
                                        compress_module comp_v_181 (
                                            .x(result[0][181]),
                                            .d(4),
                                            .result(comp_v[0][181])
                                        );
                                        
                                        compress_module comp_v_182 (
                                            .x(result[0][182]),
                                            .d(4),
                                            .result(comp_v[0][182])
                                        );
                                        
                                        compress_module comp_v_183 (
                                            .x(result[0][183]),
                                            .d(4),
                                            .result(comp_v[0][183])
                                        );
                                        
                                        compress_module comp_v_184 (
                                            .x(result[0][184]),
                                            .d(4),
                                            .result(comp_v[0][184])
                                        );
                                        
                                        compress_module comp_v_185 (
                                            .x(result[0][185]),
                                            .d(4),
                                            .result(comp_v[0][185])
                                        );
                                        
                                        compress_module comp_v_186 (
                                            .x(result[0][186]),
                                            .d(4),
                                            .result(comp_v[0][186])
                                        );
                                        
                                        compress_module comp_v_187 (
                                            .x(result[0][187]),
                                            .d(4),
                                            .result(comp_v[0][187])
                                        );
                                        
                                        compress_module comp_v_188 (
                                            .x(result[0][188]),
                                            .d(4),
                                            .result(comp_v[0][188])
                                        );
                                        
                                        compress_module comp_v_189 (
                                            .x(result[0][189]),
                                            .d(4),
                                            .result(comp_v[0][189])
                                        );
                                        
                                        compress_module comp_v_190 (
                                            .x(result[0][190]),
                                            .d(4),
                                            .result(comp_v[0][190])
                                        );
                                        
                                        compress_module comp_v_191 (
                                            .x(result[0][191]),
                                            .d(4),
                                            .result(comp_v[0][191])
                                        );
                                        
                                        compress_module comp_v_192 (
                                            .x(result[0][192]),
                                            .d(4),
                                            .result(comp_v[0][192])
                                        );
                                        
                                        compress_module comp_v_193 (
                                            .x(result[0][193]),
                                            .d(4),
                                            .result(comp_v[0][193])
                                        );
                                        
                                        compress_module comp_v_194 (
                                            .x(result[0][194]),
                                            .d(4),
                                            .result(comp_v[0][194])
                                        );
                                        
                                        compress_module comp_v_195 (
                                            .x(result[0][195]),
                                            .d(4),
                                            .result(comp_v[0][195])
                                        );
                                        
                                        compress_module comp_v_196 (
                                            .x(result[0][196]),
                                            .d(4),
                                            .result(comp_v[0][196])
                                        );
                                        
                                        compress_module comp_v_197 (
                                            .x(result[0][197]),
                                            .d(4),
                                            .result(comp_v[0][197])
                                        );
                                        
                                        compress_module comp_v_198 (
                                            .x(result[0][198]),
                                            .d(4),
                                            .result(comp_v[0][198])
                                        );
                                        
                                        compress_module comp_v_199 (
                                            .x(result[0][199]),
                                            .d(4),
                                            .result(comp_v[0][199])
                                        );
                                        
                                        compress_module comp_v_200 (
                                            .x(result[0][200]),
                                            .d(4),
                                            .result(comp_v[0][200])
                                        );
                                        
                                        compress_module comp_v_201 (
                                            .x(result[0][201]),
                                            .d(4),
                                            .result(comp_v[0][201])
                                        );
                                        
                                        compress_module comp_v_202 (
                                            .x(result[0][202]),
                                            .d(4),
                                            .result(comp_v[0][202])
                                        );
                                        
                                        compress_module comp_v_203 (
                                            .x(result[0][203]),
                                            .d(4),
                                            .result(comp_v[0][203])
                                        );
                                        
                                        compress_module comp_v_204 (
                                            .x(result[0][204]),
                                            .d(4),
                                            .result(comp_v[0][204])
                                        );
                                        
                                        compress_module comp_v_205 (
                                            .x(result[0][205]),
                                            .d(4),
                                            .result(comp_v[0][205])
                                        );
                                        
                                        compress_module comp_v_206 (
                                            .x(result[0][206]),
                                            .d(4),
                                            .result(comp_v[0][206])
                                        );
                                        
                                        compress_module comp_v_207 (
                                            .x(result[0][207]),
                                            .d(4),
                                            .result(comp_v[0][207])
                                        );
                                        
                                        compress_module comp_v_208 (
                                            .x(result[0][208]),
                                            .d(4),
                                            .result(comp_v[0][208])
                                        );
                                        
                                        compress_module comp_v_209 (
                                            .x(result[0][209]),
                                            .d(4),
                                            .result(comp_v[0][209])
                                        );
                                        
                                        compress_module comp_v_210 (
                                            .x(result[0][210]),
                                            .d(4),
                                            .result(comp_v[0][210])
                                        );
                                        
                                        compress_module comp_v_211 (
                                            .x(result[0][211]),
                                            .d(4),
                                            .result(comp_v[0][211])
                                        );
                                        
                                        compress_module comp_v_212 (
                                            .x(result[0][212]),
                                            .d(4),
                                            .result(comp_v[0][212])
                                        );
                                        
                                        compress_module comp_v_213 (
                                            .x(result[0][213]),
                                            .d(4),
                                            .result(comp_v[0][213])
                                        );
                                        
                                        compress_module comp_v_214 (
                                            .x(result[0][214]),
                                            .d(4),
                                            .result(comp_v[0][214])
                                        );
                                        
                                        compress_module comp_v_215 (
                                            .x(result[0][215]),
                                            .d(4),
                                            .result(comp_v[0][215])
                                        );
                                        
                                        compress_module comp_v_216 (
                                            .x(result[0][216]),
                                            .d(4),
                                            .result(comp_v[0][216])
                                        );
                                        
                                        compress_module comp_v_217 (
                                            .x(result[0][217]),
                                            .d(4),
                                            .result(comp_v[0][217])
                                        );
                                        
                                        compress_module comp_v_218 (
                                            .x(result[0][218]),
                                            .d(4),
                                            .result(comp_v[0][218])
                                        );
                                        
                                        compress_module comp_v_219 (
                                            .x(result[0][219]),
                                            .d(4),
                                            .result(comp_v[0][219])
                                        );
                                        
                                        compress_module comp_v_220 (
                                            .x(result[0][220]),
                                            .d(4),
                                            .result(comp_v[0][220])
                                        );
                                        
                                        compress_module comp_v_221 (
                                            .x(result[0][221]),
                                            .d(4),
                                            .result(comp_v[0][221])
                                        );
                                        
                                        compress_module comp_v_222 (
                                            .x(result[0][222]),
                                            .d(4),
                                            .result(comp_v[0][222])
                                        );
                                        
                                        compress_module comp_v_223 (
                                            .x(result[0][223]),
                                            .d(4),
                                            .result(comp_v[0][223])
                                        );
                                        
                                        compress_module comp_v_224 (
                                            .x(result[0][224]),
                                            .d(4),
                                            .result(comp_v[0][224])
                                        );
                                        
                                        compress_module comp_v_225 (
                                            .x(result[0][225]),
                                            .d(4),
                                            .result(comp_v[0][225])
                                        );
                                        
                                        compress_module comp_v_226 (
                                            .x(result[0][226]),
                                            .d(4),
                                            .result(comp_v[0][226])
                                        );
                                        
                                        compress_module comp_v_227 (
                                            .x(result[0][227]),
                                            .d(4),
                                            .result(comp_v[0][227])
                                        );
                                        
                                        compress_module comp_v_228 (
                                            .x(result[0][228]),
                                            .d(4),
                                            .result(comp_v[0][228])
                                        );
                                        
                                        compress_module comp_v_229 (
                                            .x(result[0][229]),
                                            .d(4),
                                            .result(comp_v[0][229])
                                        );
                                        
                                        compress_module comp_v_230 (
                                            .x(result[0][230]),
                                            .d(4),
                                            .result(comp_v[0][230])
                                        );
                                        
                                        compress_module comp_v_231 (
                                            .x(result[0][231]),
                                            .d(4),
                                            .result(comp_v[0][231])
                                        );
                                        
                                        compress_module comp_v_232 (
                                            .x(result[0][232]),
                                            .d(4),
                                            .result(comp_v[0][232])
                                        );
                                        
                                        compress_module comp_v_233 (
                                            .x(result[0][233]),
                                            .d(4),
                                            .result(comp_v[0][233])
                                        );
                                        
                                        compress_module comp_v_234 (
                                            .x(result[0][234]),
                                            .d(4),
                                            .result(comp_v[0][234])
                                        );
                                        
                                        compress_module comp_v_235 (
                                            .x(result[0][235]),
                                            .d(4),
                                            .result(comp_v[0][235])
                                        );
                                        
                                        compress_module comp_v_236 (
                                            .x(result[0][236]),
                                            .d(4),
                                            .result(comp_v[0][236])
                                        );
                                        
                                        compress_module comp_v_237 (
                                            .x(result[0][237]),
                                            .d(4),
                                            .result(comp_v[0][237])
                                        );
                                        
                                        compress_module comp_v_238 (
                                            .x(result[0][238]),
                                            .d(4),
                                            .result(comp_v[0][238])
                                        );
                                        
                                        compress_module comp_v_239 (
                                            .x(result[0][239]),
                                            .d(4),
                                            .result(comp_v[0][239])
                                        );
                                        
                                        compress_module comp_v_240 (
                                            .x(result[0][240]),
                                            .d(4),
                                            .result(comp_v[0][240])
                                        );
                                        
                                        compress_module comp_v_241 (
                                            .x(result[0][241]),
                                            .d(4),
                                            .result(comp_v[0][241])
                                        );
                                        
                                        compress_module comp_v_242 (
                                            .x(result[0][242]),
                                            .d(4),
                                            .result(comp_v[0][242])
                                        );
                                        
                                        compress_module comp_v_243 (
                                            .x(result[0][243]),
                                            .d(4),
                                            .result(comp_v[0][243])
                                        );
                                        
                                        compress_module comp_v_244 (
                                            .x(result[0][244]),
                                            .d(4),
                                            .result(comp_v[0][244])
                                        );
                                        
                                        compress_module comp_v_245 (
                                            .x(result[0][245]),
                                            .d(4),
                                            .result(comp_v[0][245])
                                        );
                                        
                                        compress_module comp_v_246 (
                                            .x(result[0][246]),
                                            .d(4),
                                            .result(comp_v[0][246])
                                        );
                                        
                                        compress_module comp_v_247 (
                                            .x(result[0][247]),
                                            .d(4),
                                            .result(comp_v[0][247])
                                        );
                                        
                                        compress_module comp_v_248 (
                                            .x(result[0][248]),
                                            .d(4),
                                            .result(comp_v[0][248])
                                        );
                                        
                                        compress_module comp_v_249 (
                                            .x(result[0][249]),
                                            .d(4),
                                            .result(comp_v[0][249])
                                        );
                                        
                                        compress_module comp_v_250 (
                                            .x(result[0][250]),
                                            .d(4),
                                            .result(comp_v[0][250])
                                        );
                                        
                                        compress_module comp_v_251 (
                                            .x(result[0][251]),
                                            .d(4),
                                            .result(comp_v[0][251])
                                        );
                                        
                                        compress_module comp_v_252 (
                                            .x(result[0][252]),
                                            .d(4),
                                            .result(comp_v[0][252])
                                        );
                                        
                                        compress_module comp_v_253 (
                                            .x(result[0][253]),
                                            .d(4),
                                            .result(comp_v[0][253])
                                        );
                                        
                                        compress_module comp_v_254 (
                                            .x(result[0][254]),
                                            .d(4),
                                            .result(comp_v[0][254])
                                        );
                                        
                                        compress_module comp_v_255 (
                                            .x(result[0][255]),
                                            .d(4),
                                            .result(comp_v[0][255])
                                        );
                                        
                                        compress_module comp_v_256 (
                                            .x(result[1][0]),
                                            .d(4),
                                            .result(comp_v[1][0])
                                        );
                                        
                                        compress_module comp_v_257 (
                                            .x(result[1][1]),
                                            .d(4),
                                            .result(comp_v[1][1])
                                        );
                                        
                                        compress_module comp_v_258 (
                                            .x(result[1][2]),
                                            .d(4),
                                            .result(comp_v[1][2])
                                        );
                                        
                                        compress_module comp_v_259 (
                                            .x(result[1][3]),
                                            .d(4),
                                            .result(comp_v[1][3])
                                        );
                                        
                                        compress_module comp_v_260 (
                                            .x(result[1][4]),
                                            .d(4),
                                            .result(comp_v[1][4])
                                        );
                                        
                                        compress_module comp_v_261 (
                                            .x(result[1][5]),
                                            .d(4),
                                            .result(comp_v[1][5])
                                        );
                                        
                                        compress_module comp_v_262 (
                                            .x(result[1][6]),
                                            .d(4),
                                            .result(comp_v[1][6])
                                        );
                                        
                                        compress_module comp_v_263 (
                                            .x(result[1][7]),
                                            .d(4),
                                            .result(comp_v[1][7])
                                        );
                                        
                                        compress_module comp_v_264 (
                                            .x(result[1][8]),
                                            .d(4),
                                            .result(comp_v[1][8])
                                        );
                                        
                                        compress_module comp_v_265 (
                                            .x(result[1][9]),
                                            .d(4),
                                            .result(comp_v[1][9])
                                        );
                                        
                                        compress_module comp_v_266 (
                                            .x(result[1][10]),
                                            .d(4),
                                            .result(comp_v[1][10])
                                        );
                                        
                                        compress_module comp_v_267 (
                                            .x(result[1][11]),
                                            .d(4),
                                            .result(comp_v[1][11])
                                        );
                                        
                                        compress_module comp_v_268 (
                                            .x(result[1][12]),
                                            .d(4),
                                            .result(comp_v[1][12])
                                        );
                                        
                                        compress_module comp_v_269 (
                                            .x(result[1][13]),
                                            .d(4),
                                            .result(comp_v[1][13])
                                        );
                                        
                                        compress_module comp_v_270 (
                                            .x(result[1][14]),
                                            .d(4),
                                            .result(comp_v[1][14])
                                        );
                                        
                                        compress_module comp_v_271 (
                                            .x(result[1][15]),
                                            .d(4),
                                            .result(comp_v[1][15])
                                        );
                                        
                                        compress_module comp_v_272 (
                                            .x(result[1][16]),
                                            .d(4),
                                            .result(comp_v[1][16])
                                        );
                                        
                                        compress_module comp_v_273 (
                                            .x(result[1][17]),
                                            .d(4),
                                            .result(comp_v[1][17])
                                        );
                                        
                                        compress_module comp_v_274 (
                                            .x(result[1][18]),
                                            .d(4),
                                            .result(comp_v[1][18])
                                        );
                                        
                                        compress_module comp_v_275 (
                                            .x(result[1][19]),
                                            .d(4),
                                            .result(comp_v[1][19])
                                        );
                                        
                                        compress_module comp_v_276 (
                                            .x(result[1][20]),
                                            .d(4),
                                            .result(comp_v[1][20])
                                        );
                                        
                                        compress_module comp_v_277 (
                                            .x(result[1][21]),
                                            .d(4),
                                            .result(comp_v[1][21])
                                        );
                                        
                                        compress_module comp_v_278 (
                                            .x(result[1][22]),
                                            .d(4),
                                            .result(comp_v[1][22])
                                        );
                                        
                                        compress_module comp_v_279 (
                                            .x(result[1][23]),
                                            .d(4),
                                            .result(comp_v[1][23])
                                        );
                                        
                                        compress_module comp_v_280 (
                                            .x(result[1][24]),
                                            .d(4),
                                            .result(comp_v[1][24])
                                        );
                                        
                                        compress_module comp_v_281 (
                                            .x(result[1][25]),
                                            .d(4),
                                            .result(comp_v[1][25])
                                        );
                                        
                                        compress_module comp_v_282 (
                                            .x(result[1][26]),
                                            .d(4),
                                            .result(comp_v[1][26])
                                        );
                                        
                                        compress_module comp_v_283 (
                                            .x(result[1][27]),
                                            .d(4),
                                            .result(comp_v[1][27])
                                        );
                                        
                                        compress_module comp_v_284 (
                                            .x(result[1][28]),
                                            .d(4),
                                            .result(comp_v[1][28])
                                        );
                                        
                                        compress_module comp_v_285 (
                                            .x(result[1][29]),
                                            .d(4),
                                            .result(comp_v[1][29])
                                        );
                                        
                                        compress_module comp_v_286 (
                                            .x(result[1][30]),
                                            .d(4),
                                            .result(comp_v[1][30])
                                        );
                                        
                                        compress_module comp_v_287 (
                                            .x(result[1][31]),
                                            .d(4),
                                            .result(comp_v[1][31])
                                        );
                                        
                                        compress_module comp_v_288 (
                                            .x(result[1][32]),
                                            .d(4),
                                            .result(comp_v[1][32])
                                        );
                                        
                                        compress_module comp_v_289 (
                                            .x(result[1][33]),
                                            .d(4),
                                            .result(comp_v[1][33])
                                        );
                                        
                                        compress_module comp_v_290 (
                                            .x(result[1][34]),
                                            .d(4),
                                            .result(comp_v[1][34])
                                        );
                                        
                                        compress_module comp_v_291 (
                                            .x(result[1][35]),
                                            .d(4),
                                            .result(comp_v[1][35])
                                        );
                                        
                                        compress_module comp_v_292 (
                                            .x(result[1][36]),
                                            .d(4),
                                            .result(comp_v[1][36])
                                        );
                                        
                                        compress_module comp_v_293 (
                                            .x(result[1][37]),
                                            .d(4),
                                            .result(comp_v[1][37])
                                        );
                                        
                                        compress_module comp_v_294 (
                                            .x(result[1][38]),
                                            .d(4),
                                            .result(comp_v[1][38])
                                        );
                                        
                                        compress_module comp_v_295 (
                                            .x(result[1][39]),
                                            .d(4),
                                            .result(comp_v[1][39])
                                        );
                                        
                                        compress_module comp_v_296 (
                                            .x(result[1][40]),
                                            .d(4),
                                            .result(comp_v[1][40])
                                        );
                                        
                                        compress_module comp_v_297 (
                                            .x(result[1][41]),
                                            .d(4),
                                            .result(comp_v[1][41])
                                        );
                                        
                                        compress_module comp_v_298 (
                                            .x(result[1][42]),
                                            .d(4),
                                            .result(comp_v[1][42])
                                        );
                                        
                                        compress_module comp_v_299 (
                                            .x(result[1][43]),
                                            .d(4),
                                            .result(comp_v[1][43])
                                        );
                                        
                                        compress_module comp_v_300 (
                                            .x(result[1][44]),
                                            .d(4),
                                            .result(comp_v[1][44])
                                        );
                                        
                                        compress_module comp_v_301 (
                                            .x(result[1][45]),
                                            .d(4),
                                            .result(comp_v[1][45])
                                        );
                                        
                                        compress_module comp_v_302 (
                                            .x(result[1][46]),
                                            .d(4),
                                            .result(comp_v[1][46])
                                        );
                                        
                                        compress_module comp_v_303 (
                                            .x(result[1][47]),
                                            .d(4),
                                            .result(comp_v[1][47])
                                        );
                                        
                                        compress_module comp_v_304 (
                                            .x(result[1][48]),
                                            .d(4),
                                            .result(comp_v[1][48])
                                        );
                                        
                                        compress_module comp_v_305 (
                                            .x(result[1][49]),
                                            .d(4),
                                            .result(comp_v[1][49])
                                        );
                                        
                                        compress_module comp_v_306 (
                                            .x(result[1][50]),
                                            .d(4),
                                            .result(comp_v[1][50])
                                        );
                                        
                                        compress_module comp_v_307 (
                                            .x(result[1][51]),
                                            .d(4),
                                            .result(comp_v[1][51])
                                        );
                                        
                                        compress_module comp_v_308 (
                                            .x(result[1][52]),
                                            .d(4),
                                            .result(comp_v[1][52])
                                        );
                                        
                                        compress_module comp_v_309 (
                                            .x(result[1][53]),
                                            .d(4),
                                            .result(comp_v[1][53])
                                        );
                                        
                                        compress_module comp_v_310 (
                                            .x(result[1][54]),
                                            .d(4),
                                            .result(comp_v[1][54])
                                        );
                                        
                                        compress_module comp_v_311 (
                                            .x(result[1][55]),
                                            .d(4),
                                            .result(comp_v[1][55])
                                        );
                                        
                                        compress_module comp_v_312 (
                                            .x(result[1][56]),
                                            .d(4),
                                            .result(comp_v[1][56])
                                        );
                                        
                                        compress_module comp_v_313 (
                                            .x(result[1][57]),
                                            .d(4),
                                            .result(comp_v[1][57])
                                        );
                                        
                                        compress_module comp_v_314 (
                                            .x(result[1][58]),
                                            .d(4),
                                            .result(comp_v[1][58])
                                        );
                                        
                                        compress_module comp_v_315 (
                                            .x(result[1][59]),
                                            .d(4),
                                            .result(comp_v[1][59])
                                        );
                                        
                                        compress_module comp_v_316 (
                                            .x(result[1][60]),
                                            .d(4),
                                            .result(comp_v[1][60])
                                        );
                                        
                                        compress_module comp_v_317 (
                                            .x(result[1][61]),
                                            .d(4),
                                            .result(comp_v[1][61])
                                        );
                                        
                                        compress_module comp_v_318 (
                                            .x(result[1][62]),
                                            .d(4),
                                            .result(comp_v[1][62])
                                        );
                                        
                                        compress_module comp_v_319 (
                                            .x(result[1][63]),
                                            .d(4),
                                            .result(comp_v[1][63])
                                        );
                                        
                                        compress_module comp_v_320 (
                                            .x(result[1][64]),
                                            .d(4),
                                            .result(comp_v[1][64])
                                        );
                                        
                                        compress_module comp_v_321 (
                                            .x(result[1][65]),
                                            .d(4),
                                            .result(comp_v[1][65])
                                        );
                                        
                                        compress_module comp_v_322 (
                                            .x(result[1][66]),
                                            .d(4),
                                            .result(comp_v[1][66])
                                        );
                                        
                                        compress_module comp_v_323 (
                                            .x(result[1][67]),
                                            .d(4),
                                            .result(comp_v[1][67])
                                        );
                                        
                                        compress_module comp_v_324 (
                                            .x(result[1][68]),
                                            .d(4),
                                            .result(comp_v[1][68])
                                        );
                                        
                                        compress_module comp_v_325 (
                                            .x(result[1][69]),
                                            .d(4),
                                            .result(comp_v[1][69])
                                        );
                                        
                                        compress_module comp_v_326 (
                                            .x(result[1][70]),
                                            .d(4),
                                            .result(comp_v[1][70])
                                        );
                                        
                                        compress_module comp_v_327 (
                                            .x(result[1][71]),
                                            .d(4),
                                            .result(comp_v[1][71])
                                        );
                                        
                                        compress_module comp_v_328 (
                                            .x(result[1][72]),
                                            .d(4),
                                            .result(comp_v[1][72])
                                        );
                                        
                                        compress_module comp_v_329 (
                                            .x(result[1][73]),
                                            .d(4),
                                            .result(comp_v[1][73])
                                        );
                                        
                                        compress_module comp_v_330 (
                                            .x(result[1][74]),
                                            .d(4),
                                            .result(comp_v[1][74])
                                        );
                                        
                                        compress_module comp_v_331 (
                                            .x(result[1][75]),
                                            .d(4),
                                            .result(comp_v[1][75])
                                        );
                                        
                                        compress_module comp_v_332 (
                                            .x(result[1][76]),
                                            .d(4),
                                            .result(comp_v[1][76])
                                        );
                                        
                                        compress_module comp_v_333 (
                                            .x(result[1][77]),
                                            .d(4),
                                            .result(comp_v[1][77])
                                        );
                                        
                                        compress_module comp_v_334 (
                                            .x(result[1][78]),
                                            .d(4),
                                            .result(comp_v[1][78])
                                        );
                                        
                                        compress_module comp_v_335 (
                                            .x(result[1][79]),
                                            .d(4),
                                            .result(comp_v[1][79])
                                        );
                                        
                                        compress_module comp_v_336 (
                                            .x(result[1][80]),
                                            .d(4),
                                            .result(comp_v[1][80])
                                        );
                                        
                                        compress_module comp_v_337 (
                                            .x(result[1][81]),
                                            .d(4),
                                            .result(comp_v[1][81])
                                        );
                                        
                                        compress_module comp_v_338 (
                                            .x(result[1][82]),
                                            .d(4),
                                            .result(comp_v[1][82])
                                        );
                                        
                                        compress_module comp_v_339 (
                                            .x(result[1][83]),
                                            .d(4),
                                            .result(comp_v[1][83])
                                        );
                                        
                                        compress_module comp_v_340 (
                                            .x(result[1][84]),
                                            .d(4),
                                            .result(comp_v[1][84])
                                        );
                                        
                                        compress_module comp_v_341 (
                                            .x(result[1][85]),
                                            .d(4),
                                            .result(comp_v[1][85])
                                        );
                                        
                                        compress_module comp_v_342 (
                                            .x(result[1][86]),
                                            .d(4),
                                            .result(comp_v[1][86])
                                        );
                                        
                                        compress_module comp_v_343 (
                                            .x(result[1][87]),
                                            .d(4),
                                            .result(comp_v[1][87])
                                        );
                                        
                                        compress_module comp_v_344 (
                                            .x(result[1][88]),
                                            .d(4),
                                            .result(comp_v[1][88])
                                        );
                                        
                                        compress_module comp_v_345 (
                                            .x(result[1][89]),
                                            .d(4),
                                            .result(comp_v[1][89])
                                        );
                                        
                                        compress_module comp_v_346 (
                                            .x(result[1][90]),
                                            .d(4),
                                            .result(comp_v[1][90])
                                        );
                                        
                                        compress_module comp_v_347 (
                                            .x(result[1][91]),
                                            .d(4),
                                            .result(comp_v[1][91])
                                        );
                                        
                                        compress_module comp_v_348 (
                                            .x(result[1][92]),
                                            .d(4),
                                            .result(comp_v[1][92])
                                        );
                                        
                                        compress_module comp_v_349 (
                                            .x(result[1][93]),
                                            .d(4),
                                            .result(comp_v[1][93])
                                        );
                                        
                                        compress_module comp_v_350 (
                                            .x(result[1][94]),
                                            .d(4),
                                            .result(comp_v[1][94])
                                        );
                                        
                                        compress_module comp_v_351 (
                                            .x(result[1][95]),
                                            .d(4),
                                            .result(comp_v[1][95])
                                        );
                                        
                                        compress_module comp_v_352 (
                                            .x(result[1][96]),
                                            .d(4),
                                            .result(comp_v[1][96])
                                        );
                                        
                                        compress_module comp_v_353 (
                                            .x(result[1][97]),
                                            .d(4),
                                            .result(comp_v[1][97])
                                        );
                                        
                                        compress_module comp_v_354 (
                                            .x(result[1][98]),
                                            .d(4),
                                            .result(comp_v[1][98])
                                        );
                                        
                                        compress_module comp_v_355 (
                                            .x(result[1][99]),
                                            .d(4),
                                            .result(comp_v[1][99])
                                        );
                                        
                                        compress_module comp_v_356 (
                                            .x(result[1][100]),
                                            .d(4),
                                            .result(comp_v[1][100])
                                        );
                                        
                                        compress_module comp_v_357 (
                                            .x(result[1][101]),
                                            .d(4),
                                            .result(comp_v[1][101])
                                        );
                                        
                                        compress_module comp_v_358 (
                                            .x(result[1][102]),
                                            .d(4),
                                            .result(comp_v[1][102])
                                        );
                                        
                                        compress_module comp_v_359 (
                                            .x(result[1][103]),
                                            .d(4),
                                            .result(comp_v[1][103])
                                        );
                                        
                                        compress_module comp_v_360 (
                                            .x(result[1][104]),
                                            .d(4),
                                            .result(comp_v[1][104])
                                        );
                                        
                                        compress_module comp_v_361 (
                                            .x(result[1][105]),
                                            .d(4),
                                            .result(comp_v[1][105])
                                        );
                                        
                                        compress_module comp_v_362 (
                                            .x(result[1][106]),
                                            .d(4),
                                            .result(comp_v[1][106])
                                        );
                                        
                                        compress_module comp_v_363 (
                                            .x(result[1][107]),
                                            .d(4),
                                            .result(comp_v[1][107])
                                        );
                                        
                                        compress_module comp_v_364 (
                                            .x(result[1][108]),
                                            .d(4),
                                            .result(comp_v[1][108])
                                        );
                                        
                                        compress_module comp_v_365 (
                                            .x(result[1][109]),
                                            .d(4),
                                            .result(comp_v[1][109])
                                        );
                                        
                                        compress_module comp_v_366 (
                                            .x(result[1][110]),
                                            .d(4),
                                            .result(comp_v[1][110])
                                        );
                                        
                                        compress_module comp_v_367 (
                                            .x(result[1][111]),
                                            .d(4),
                                            .result(comp_v[1][111])
                                        );
                                        
                                        compress_module comp_v_368 (
                                            .x(result[1][112]),
                                            .d(4),
                                            .result(comp_v[1][112])
                                        );
                                        
                                        compress_module comp_v_369 (
                                            .x(result[1][113]),
                                            .d(4),
                                            .result(comp_v[1][113])
                                        );
                                        
                                        compress_module comp_v_370 (
                                            .x(result[1][114]),
                                            .d(4),
                                            .result(comp_v[1][114])
                                        );
                                        
                                        compress_module comp_v_371 (
                                            .x(result[1][115]),
                                            .d(4),
                                            .result(comp_v[1][115])
                                        );
                                        
                                        compress_module comp_v_372 (
                                            .x(result[1][116]),
                                            .d(4),
                                            .result(comp_v[1][116])
                                        );
                                        
                                        compress_module comp_v_373 (
                                            .x(result[1][117]),
                                            .d(4),
                                            .result(comp_v[1][117])
                                        );
                                        
                                        compress_module comp_v_374 (
                                            .x(result[1][118]),
                                            .d(4),
                                            .result(comp_v[1][118])
                                        );
                                        
                                        compress_module comp_v_375 (
                                            .x(result[1][119]),
                                            .d(4),
                                            .result(comp_v[1][119])
                                        );
                                        
                                        compress_module comp_v_376 (
                                            .x(result[1][120]),
                                            .d(4),
                                            .result(comp_v[1][120])
                                        );
                                        
                                        compress_module comp_v_377 (
                                            .x(result[1][121]),
                                            .d(4),
                                            .result(comp_v[1][121])
                                        );
                                        
                                        compress_module comp_v_378 (
                                            .x(result[1][122]),
                                            .d(4),
                                            .result(comp_v[1][122])
                                        );
                                        
                                        compress_module comp_v_379 (
                                            .x(result[1][123]),
                                            .d(4),
                                            .result(comp_v[1][123])
                                        );
                                        
                                        compress_module comp_v_380 (
                                            .x(result[1][124]),
                                            .d(4),
                                            .result(comp_v[1][124])
                                        );
                                        
                                        compress_module comp_v_381 (
                                            .x(result[1][125]),
                                            .d(4),
                                            .result(comp_v[1][125])
                                        );
                                        
                                        compress_module comp_v_382 (
                                            .x(result[1][126]),
                                            .d(4),
                                            .result(comp_v[1][126])
                                        );
                                        
                                        compress_module comp_v_383 (
                                            .x(result[1][127]),
                                            .d(4),
                                            .result(comp_v[1][127])
                                        );
                                        
                                        compress_module comp_v_384 (
                                            .x(result[1][128]),
                                            .d(4),
                                            .result(comp_v[1][128])
                                        );
                                        
                                        compress_module comp_v_385 (
                                            .x(result[1][129]),
                                            .d(4),
                                            .result(comp_v[1][129])
                                        );
                                        
                                        compress_module comp_v_386 (
                                            .x(result[1][130]),
                                            .d(4),
                                            .result(comp_v[1][130])
                                        );
                                        
                                        compress_module comp_v_387 (
                                            .x(result[1][131]),
                                            .d(4),
                                            .result(comp_v[1][131])
                                        );
                                        
                                        compress_module comp_v_388 (
                                            .x(result[1][132]),
                                            .d(4),
                                            .result(comp_v[1][132])
                                        );
                                        
                                        compress_module comp_v_389 (
                                            .x(result[1][133]),
                                            .d(4),
                                            .result(comp_v[1][133])
                                        );
                                        
                                        compress_module comp_v_390 (
                                            .x(result[1][134]),
                                            .d(4),
                                            .result(comp_v[1][134])
                                        );
                                        
                                        compress_module comp_v_391 (
                                            .x(result[1][135]),
                                            .d(4),
                                            .result(comp_v[1][135])
                                        );
                                        
                                        compress_module comp_v_392 (
                                            .x(result[1][136]),
                                            .d(4),
                                            .result(comp_v[1][136])
                                        );
                                        
                                        compress_module comp_v_393 (
                                            .x(result[1][137]),
                                            .d(4),
                                            .result(comp_v[1][137])
                                        );
                                        
                                        compress_module comp_v_394 (
                                            .x(result[1][138]),
                                            .d(4),
                                            .result(comp_v[1][138])
                                        );
                                        
                                        compress_module comp_v_395 (
                                            .x(result[1][139]),
                                            .d(4),
                                            .result(comp_v[1][139])
                                        );
                                        
                                        compress_module comp_v_396 (
                                            .x(result[1][140]),
                                            .d(4),
                                            .result(comp_v[1][140])
                                        );
                                        
                                        compress_module comp_v_397 (
                                            .x(result[1][141]),
                                            .d(4),
                                            .result(comp_v[1][141])
                                        );
                                        
                                        compress_module comp_v_398 (
                                            .x(result[1][142]),
                                            .d(4),
                                            .result(comp_v[1][142])
                                        );
                                        
                                        compress_module comp_v_399 (
                                            .x(result[1][143]),
                                            .d(4),
                                            .result(comp_v[1][143])
                                        );
                                        
                                        compress_module comp_v_400 (
                                            .x(result[1][144]),
                                            .d(4),
                                            .result(comp_v[1][144])
                                        );
                                        
                                        compress_module comp_v_401 (
                                            .x(result[1][145]),
                                            .d(4),
                                            .result(comp_v[1][145])
                                        );
                                        
                                        compress_module comp_v_402 (
                                            .x(result[1][146]),
                                            .d(4),
                                            .result(comp_v[1][146])
                                        );
                                        
                                        compress_module comp_v_403 (
                                            .x(result[1][147]),
                                            .d(4),
                                            .result(comp_v[1][147])
                                        );
                                        
                                        compress_module comp_v_404 (
                                            .x(result[1][148]),
                                            .d(4),
                                            .result(comp_v[1][148])
                                        );
                                        
                                        compress_module comp_v_405 (
                                            .x(result[1][149]),
                                            .d(4),
                                            .result(comp_v[1][149])
                                        );
                                        
                                        compress_module comp_v_406 (
                                            .x(result[1][150]),
                                            .d(4),
                                            .result(comp_v[1][150])
                                        );
                                        
                                        compress_module comp_v_407 (
                                            .x(result[1][151]),
                                            .d(4),
                                            .result(comp_v[1][151])
                                        );
                                        
                                        compress_module comp_v_408 (
                                            .x(result[1][152]),
                                            .d(4),
                                            .result(comp_v[1][152])
                                        );
                                        
                                        compress_module comp_v_409 (
                                            .x(result[1][153]),
                                            .d(4),
                                            .result(comp_v[1][153])
                                        );
                                        
                                        compress_module comp_v_410 (
                                            .x(result[1][154]),
                                            .d(4),
                                            .result(comp_v[1][154])
                                        );
                                        
                                        compress_module comp_v_411 (
                                            .x(result[1][155]),
                                            .d(4),
                                            .result(comp_v[1][155])
                                        );
                                        
                                        compress_module comp_v_412 (
                                            .x(result[1][156]),
                                            .d(4),
                                            .result(comp_v[1][156])
                                        );
                                        
                                        compress_module comp_v_413 (
                                            .x(result[1][157]),
                                            .d(4),
                                            .result(comp_v[1][157])
                                        );
                                        
                                        compress_module comp_v_414 (
                                            .x(result[1][158]),
                                            .d(4),
                                            .result(comp_v[1][158])
                                        );
                                        
                                        compress_module comp_v_415 (
                                            .x(result[1][159]),
                                            .d(4),
                                            .result(comp_v[1][159])
                                        );
                                        
                                        compress_module comp_v_416 (
                                            .x(result[1][160]),
                                            .d(4),
                                            .result(comp_v[1][160])
                                        );
                                        
                                        compress_module comp_v_417 (
                                            .x(result[1][161]),
                                            .d(4),
                                            .result(comp_v[1][161])
                                        );
                                        
                                        compress_module comp_v_418 (
                                            .x(result[1][162]),
                                            .d(4),
                                            .result(comp_v[1][162])
                                        );
                                        
                                        compress_module comp_v_419 (
                                            .x(result[1][163]),
                                            .d(4),
                                            .result(comp_v[1][163])
                                        );
                                        
                                        compress_module comp_v_420 (
                                            .x(result[1][164]),
                                            .d(4),
                                            .result(comp_v[1][164])
                                        );
                                        
                                        compress_module comp_v_421 (
                                            .x(result[1][165]),
                                            .d(4),
                                            .result(comp_v[1][165])
                                        );
                                        
                                        compress_module comp_v_422 (
                                            .x(result[1][166]),
                                            .d(4),
                                            .result(comp_v[1][166])
                                        );
                                        
                                        compress_module comp_v_423 (
                                            .x(result[1][167]),
                                            .d(4),
                                            .result(comp_v[1][167])
                                        );
                                        
                                        compress_module comp_v_424 (
                                            .x(result[1][168]),
                                            .d(4),
                                            .result(comp_v[1][168])
                                        );
                                        
                                        compress_module comp_v_425 (
                                            .x(result[1][169]),
                                            .d(4),
                                            .result(comp_v[1][169])
                                        );
                                        
                                        compress_module comp_v_426 (
                                            .x(result[1][170]),
                                            .d(4),
                                            .result(comp_v[1][170])
                                        );
                                        
                                        compress_module comp_v_427 (
                                            .x(result[1][171]),
                                            .d(4),
                                            .result(comp_v[1][171])
                                        );
                                        
                                        compress_module comp_v_428 (
                                            .x(result[1][172]),
                                            .d(4),
                                            .result(comp_v[1][172])
                                        );
                                        
                                        compress_module comp_v_429 (
                                            .x(result[1][173]),
                                            .d(4),
                                            .result(comp_v[1][173])
                                        );
                                        
                                        compress_module comp_v_430 (
                                            .x(result[1][174]),
                                            .d(4),
                                            .result(comp_v[1][174])
                                        );
                                        
                                        compress_module comp_v_431 (
                                            .x(result[1][175]),
                                            .d(4),
                                            .result(comp_v[1][175])
                                        );
                                        
                                        compress_module comp_v_432 (
                                            .x(result[1][176]),
                                            .d(4),
                                            .result(comp_v[1][176])
                                        );
                                        
                                        compress_module comp_v_433 (
                                            .x(result[1][177]),
                                            .d(4),
                                            .result(comp_v[1][177])
                                        );
                                        
                                        compress_module comp_v_434 (
                                            .x(result[1][178]),
                                            .d(4),
                                            .result(comp_v[1][178])
                                        );
                                        
                                        compress_module comp_v_435 (
                                            .x(result[1][179]),
                                            .d(4),
                                            .result(comp_v[1][179])
                                        );
                                        
                                        compress_module comp_v_436 (
                                            .x(result[1][180]),
                                            .d(4),
                                            .result(comp_v[1][180])
                                        );
                                        
                                        compress_module comp_v_437 (
                                            .x(result[1][181]),
                                            .d(4),
                                            .result(comp_v[1][181])
                                        );
                                        
                                        compress_module comp_v_438 (
                                            .x(result[1][182]),
                                            .d(4),
                                            .result(comp_v[1][182])
                                        );
                                        
                                        compress_module comp_v_439 (
                                            .x(result[1][183]),
                                            .d(4),
                                            .result(comp_v[1][183])
                                        );
                                        
                                        compress_module comp_v_440 (
                                            .x(result[1][184]),
                                            .d(4),
                                            .result(comp_v[1][184])
                                        );
                                        
                                        compress_module comp_v_441 (
                                            .x(result[1][185]),
                                            .d(4),
                                            .result(comp_v[1][185])
                                        );
                                        
                                        compress_module comp_v_442 (
                                            .x(result[1][186]),
                                            .d(4),
                                            .result(comp_v[1][186])
                                        );
                                        
                                        compress_module comp_v_443 (
                                            .x(result[1][187]),
                                            .d(4),
                                            .result(comp_v[1][187])
                                        );
                                        
                                        compress_module comp_v_444 (
                                            .x(result[1][188]),
                                            .d(4),
                                            .result(comp_v[1][188])
                                        );
                                        
                                        compress_module comp_v_445 (
                                            .x(result[1][189]),
                                            .d(4),
                                            .result(comp_v[1][189])
                                        );
                                        
                                        compress_module comp_v_446 (
                                            .x(result[1][190]),
                                            .d(4),
                                            .result(comp_v[1][190])
                                        );
                                        
                                        compress_module comp_v_447 (
                                            .x(result[1][191]),
                                            .d(4),
                                            .result(comp_v[1][191])
                                        );
                                        
                                        compress_module comp_v_448 (
                                            .x(result[1][192]),
                                            .d(4),
                                            .result(comp_v[1][192])
                                        );
                                        
                                        compress_module comp_v_449 (
                                            .x(result[1][193]),
                                            .d(4),
                                            .result(comp_v[1][193])
                                        );
                                        
                                        compress_module comp_v_450 (
                                            .x(result[1][194]),
                                            .d(4),
                                            .result(comp_v[1][194])
                                        );
                                        
                                        compress_module comp_v_451 (
                                            .x(result[1][195]),
                                            .d(4),
                                            .result(comp_v[1][195])
                                        );
                                        
                                        compress_module comp_v_452 (
                                            .x(result[1][196]),
                                            .d(4),
                                            .result(comp_v[1][196])
                                        );
                                        
                                        compress_module comp_v_453 (
                                            .x(result[1][197]),
                                            .d(4),
                                            .result(comp_v[1][197])
                                        );
                                        
                                        compress_module comp_v_454 (
                                            .x(result[1][198]),
                                            .d(4),
                                            .result(comp_v[1][198])
                                        );
                                        
                                        compress_module comp_v_455 (
                                            .x(result[1][199]),
                                            .d(4),
                                            .result(comp_v[1][199])
                                        );
                                        
                                        compress_module comp_v_456 (
                                            .x(result[1][200]),
                                            .d(4),
                                            .result(comp_v[1][200])
                                        );
                                        
                                        compress_module comp_v_457 (
                                            .x(result[1][201]),
                                            .d(4),
                                            .result(comp_v[1][201])
                                        );
                                        
                                        compress_module comp_v_458 (
                                            .x(result[1][202]),
                                            .d(4),
                                            .result(comp_v[1][202])
                                        );
                                        
                                        compress_module comp_v_459 (
                                            .x(result[1][203]),
                                            .d(4),
                                            .result(comp_v[1][203])
                                        );
                                        
                                        compress_module comp_v_460 (
                                            .x(result[1][204]),
                                            .d(4),
                                            .result(comp_v[1][204])
                                        );
                                        
                                        compress_module comp_v_461 (
                                            .x(result[1][205]),
                                            .d(4),
                                            .result(comp_v[1][205])
                                        );
                                        
                                        compress_module comp_v_462 (
                                            .x(result[1][206]),
                                            .d(4),
                                            .result(comp_v[1][206])
                                        );
                                        
                                        compress_module comp_v_463 (
                                            .x(result[1][207]),
                                            .d(4),
                                            .result(comp_v[1][207])
                                        );
                                        
                                        compress_module comp_v_464 (
                                            .x(result[1][208]),
                                            .d(4),
                                            .result(comp_v[1][208])
                                        );
                                        
                                        compress_module comp_v_465 (
                                            .x(result[1][209]),
                                            .d(4),
                                            .result(comp_v[1][209])
                                        );
                                        
                                        compress_module comp_v_466 (
                                            .x(result[1][210]),
                                            .d(4),
                                            .result(comp_v[1][210])
                                        );
                                        
                                        compress_module comp_v_467 (
                                            .x(result[1][211]),
                                            .d(4),
                                            .result(comp_v[1][211])
                                        );
                                        
                                        compress_module comp_v_468 (
                                            .x(result[1][212]),
                                            .d(4),
                                            .result(comp_v[1][212])
                                        );
                                        
                                        compress_module comp_v_469 (
                                            .x(result[1][213]),
                                            .d(4),
                                            .result(comp_v[1][213])
                                        );
                                        
                                        compress_module comp_v_470 (
                                            .x(result[1][214]),
                                            .d(4),
                                            .result(comp_v[1][214])
                                        );
                                        
                                        compress_module comp_v_471 (
                                            .x(result[1][215]),
                                            .d(4),
                                            .result(comp_v[1][215])
                                        );
                                        
                                        compress_module comp_v_472 (
                                            .x(result[1][216]),
                                            .d(4),
                                            .result(comp_v[1][216])
                                        );
                                        
                                        compress_module comp_v_473 (
                                            .x(result[1][217]),
                                            .d(4),
                                            .result(comp_v[1][217])
                                        );
                                        
                                        compress_module comp_v_474 (
                                            .x(result[1][218]),
                                            .d(4),
                                            .result(comp_v[1][218])
                                        );
                                        
                                        compress_module comp_v_475 (
                                            .x(result[1][219]),
                                            .d(4),
                                            .result(comp_v[1][219])
                                        );
                                        
                                        compress_module comp_v_476 (
                                            .x(result[1][220]),
                                            .d(4),
                                            .result(comp_v[1][220])
                                        );
                                        
                                        compress_module comp_v_477 (
                                            .x(result[1][221]),
                                            .d(4),
                                            .result(comp_v[1][221])
                                        );
                                        
                                        compress_module comp_v_478 (
                                            .x(result[1][222]),
                                            .d(4),
                                            .result(comp_v[1][222])
                                        );
                                        
                                        compress_module comp_v_479 (
                                            .x(result[1][223]),
                                            .d(4),
                                            .result(comp_v[1][223])
                                        );
                                        
                                        compress_module comp_v_480 (
                                            .x(result[1][224]),
                                            .d(4),
                                            .result(comp_v[1][224])
                                        );
                                        
                                        compress_module comp_v_481 (
                                            .x(result[1][225]),
                                            .d(4),
                                            .result(comp_v[1][225])
                                        );
                                        
                                        compress_module comp_v_482 (
                                            .x(result[1][226]),
                                            .d(4),
                                            .result(comp_v[1][226])
                                        );
                                        
                                        compress_module comp_v_483 (
                                            .x(result[1][227]),
                                            .d(4),
                                            .result(comp_v[1][227])
                                        );
                                        
                                        compress_module comp_v_484 (
                                            .x(result[1][228]),
                                            .d(4),
                                            .result(comp_v[1][228])
                                        );
                                        
                                        compress_module comp_v_485 (
                                            .x(result[1][229]),
                                            .d(4),
                                            .result(comp_v[1][229])
                                        );
                                        
                                        compress_module comp_v_486 (
                                            .x(result[1][230]),
                                            .d(4),
                                            .result(comp_v[1][230])
                                        );
                                        
                                        compress_module comp_v_487 (
                                            .x(result[1][231]),
                                            .d(4),
                                            .result(comp_v[1][231])
                                        );
                                        
                                        compress_module comp_v_488 (
                                            .x(result[1][232]),
                                            .d(4),
                                            .result(comp_v[1][232])
                                        );
                                        
                                        compress_module comp_v_489 (
                                            .x(result[1][233]),
                                            .d(4),
                                            .result(comp_v[1][233])
                                        );
                                        
                                        compress_module comp_v_490 (
                                            .x(result[1][234]),
                                            .d(4),
                                            .result(comp_v[1][234])
                                        );
                                        
                                        compress_module comp_v_491 (
                                            .x(result[1][235]),
                                            .d(4),
                                            .result(comp_v[1][235])
                                        );
                                        
                                        compress_module comp_v_492 (
                                            .x(result[1][236]),
                                            .d(4),
                                            .result(comp_v[1][236])
                                        );
                                        
                                        compress_module comp_v_493 (
                                            .x(result[1][237]),
                                            .d(4),
                                            .result(comp_v[1][237])
                                        );
                                        
                                        compress_module comp_v_494 (
                                            .x(result[1][238]),
                                            .d(4),
                                            .result(comp_v[1][238])
                                        );
                                        
                                        compress_module comp_v_495 (
                                            .x(result[1][239]),
                                            .d(4),
                                            .result(comp_v[1][239])
                                        );
                                        
                                        compress_module comp_v_496 (
                                            .x(result[1][240]),
                                            .d(4),
                                            .result(comp_v[1][240])
                                        );
                                        
                                        compress_module comp_v_497 (
                                            .x(result[1][241]),
                                            .d(4),
                                            .result(comp_v[1][241])
                                        );
                                        
                                        compress_module comp_v_498 (
                                            .x(result[1][242]),
                                            .d(4),
                                            .result(comp_v[1][242])
                                        );
                                        
                                        compress_module comp_v_499 (
                                            .x(result[1][243]),
                                            .d(4),
                                            .result(comp_v[1][243])
                                        );
                                        
                                        compress_module comp_v_500 (
                                            .x(result[1][244]),
                                            .d(4),
                                            .result(comp_v[1][244])
                                        );
                                        
                                        compress_module comp_v_501 (
                                            .x(result[1][245]),
                                            .d(4),
                                            .result(comp_v[1][245])
                                        );
                                        
                                        compress_module comp_v_502 (
                                            .x(result[1][246]),
                                            .d(4),
                                            .result(comp_v[1][246])
                                        );
                                        
                                        compress_module comp_v_503 (
                                            .x(result[1][247]),
                                            .d(4),
                                            .result(comp_v[1][247])
                                        );
                                        
                                        compress_module comp_v_504 (
                                            .x(result[1][248]),
                                            .d(4),
                                            .result(comp_v[1][248])
                                        );
                                        
                                        compress_module comp_v_505 (
                                            .x(result[1][249]),
                                            .d(4),
                                            .result(comp_v[1][249])
                                        );
                                        
                                        compress_module comp_v_506 (
                                            .x(result[1][250]),
                                            .d(4),
                                            .result(comp_v[1][250])
                                        );
                                        
                                        compress_module comp_v_507 (
                                            .x(result[1][251]),
                                            .d(4),
                                            .result(comp_v[1][251])
                                        );
                                        
                                        compress_module comp_v_508 (
                                            .x(result[1][252]),
                                            .d(4),
                                            .result(comp_v[1][252])
                                        );
                                        
                                        compress_module comp_v_509 (
                                            .x(result[1][253]),
                                            .d(4),
                                            .result(comp_v[1][253])
                                        );
                                        
                                        compress_module comp_v_510 (
                                            .x(result[1][254]),
                                            .d(4),
                                            .result(comp_v[1][254])
                                        );
                                        
                                        compress_module comp_v_511 (
                                            .x(result[1][255]),
                                            .d(4),
                                            .result(comp_v[1][255])
                                        );
                                        
                                        compress_module comp_v_512 (
                                            .x(result[2][0]),
                                            .d(4),
                                            .result(comp_v[2][0])
                                        );
                                        
                                        compress_module comp_v_513 (
                                            .x(result[2][1]),
                                            .d(4),
                                            .result(comp_v[2][1])
                                        );
                                        
                                        compress_module comp_v_514 (
                                            .x(result[2][2]),
                                            .d(4),
                                            .result(comp_v[2][2])
                                        );
                                        
                                        compress_module comp_v_515 (
                                            .x(result[2][3]),
                                            .d(4),
                                            .result(comp_v[2][3])
                                        );
                                        
                                        compress_module comp_v_516 (
                                            .x(result[2][4]),
                                            .d(4),
                                            .result(comp_v[2][4])
                                        );
                                        
                                        compress_module comp_v_517 (
                                            .x(result[2][5]),
                                            .d(4),
                                            .result(comp_v[2][5])
                                        );
                                        
                                        compress_module comp_v_518 (
                                            .x(result[2][6]),
                                            .d(4),
                                            .result(comp_v[2][6])
                                        );
                                        
                                        compress_module comp_v_519 (
                                            .x(result[2][7]),
                                            .d(4),
                                            .result(comp_v[2][7])
                                        );
                                        
                                        compress_module comp_v_520 (
                                            .x(result[2][8]),
                                            .d(4),
                                            .result(comp_v[2][8])
                                        );
                                        
                                        compress_module comp_v_521 (
                                            .x(result[2][9]),
                                            .d(4),
                                            .result(comp_v[2][9])
                                        );
                                        
                                        compress_module comp_v_522 (
                                            .x(result[2][10]),
                                            .d(4),
                                            .result(comp_v[2][10])
                                        );
                                        
                                        compress_module comp_v_523 (
                                            .x(result[2][11]),
                                            .d(4),
                                            .result(comp_v[2][11])
                                        );
                                        
                                        compress_module comp_v_524 (
                                            .x(result[2][12]),
                                            .d(4),
                                            .result(comp_v[2][12])
                                        );
                                        
                                        compress_module comp_v_525 (
                                            .x(result[2][13]),
                                            .d(4),
                                            .result(comp_v[2][13])
                                        );
                                        
                                        compress_module comp_v_526 (
                                            .x(result[2][14]),
                                            .d(4),
                                            .result(comp_v[2][14])
                                        );
                                        
                                        compress_module comp_v_527 (
                                            .x(result[2][15]),
                                            .d(4),
                                            .result(comp_v[2][15])
                                        );
                                        
                                        compress_module comp_v_528 (
                                            .x(result[2][16]),
                                            .d(4),
                                            .result(comp_v[2][16])
                                        );
                                        
                                        compress_module comp_v_529 (
                                            .x(result[2][17]),
                                            .d(4),
                                            .result(comp_v[2][17])
                                        );
                                        
                                        compress_module comp_v_530 (
                                            .x(result[2][18]),
                                            .d(4),
                                            .result(comp_v[2][18])
                                        );
                                        
                                        compress_module comp_v_531 (
                                            .x(result[2][19]),
                                            .d(4),
                                            .result(comp_v[2][19])
                                        );
                                        
                                        compress_module comp_v_532 (
                                            .x(result[2][20]),
                                            .d(4),
                                            .result(comp_v[2][20])
                                        );
                                        
                                        compress_module comp_v_533 (
                                            .x(result[2][21]),
                                            .d(4),
                                            .result(comp_v[2][21])
                                        );
                                        
                                        compress_module comp_v_534 (
                                            .x(result[2][22]),
                                            .d(4),
                                            .result(comp_v[2][22])
                                        );
                                        
                                        compress_module comp_v_535 (
                                            .x(result[2][23]),
                                            .d(4),
                                            .result(comp_v[2][23])
                                        );
                                        
                                        compress_module comp_v_536 (
                                            .x(result[2][24]),
                                            .d(4),
                                            .result(comp_v[2][24])
                                        );
                                        
                                        compress_module comp_v_537 (
                                            .x(result[2][25]),
                                            .d(4),
                                            .result(comp_v[2][25])
                                        );
                                        
                                        compress_module comp_v_538 (
                                            .x(result[2][26]),
                                            .d(4),
                                            .result(comp_v[2][26])
                                        );
                                        
                                        compress_module comp_v_539 (
                                            .x(result[2][27]),
                                            .d(4),
                                            .result(comp_v[2][27])
                                        );
                                        
                                        compress_module comp_v_540 (
                                            .x(result[2][28]),
                                            .d(4),
                                            .result(comp_v[2][28])
                                        );
                                        
                                        compress_module comp_v_541 (
                                            .x(result[2][29]),
                                            .d(4),
                                            .result(comp_v[2][29])
                                        );
                                        
                                        compress_module comp_v_542 (
                                            .x(result[2][30]),
                                            .d(4),
                                            .result(comp_v[2][30])
                                        );
                                        
                                        compress_module comp_v_543 (
                                            .x(result[2][31]),
                                            .d(4),
                                            .result(comp_v[2][31])
                                        );
                                        
                                        compress_module comp_v_544 (
                                            .x(result[2][32]),
                                            .d(4),
                                            .result(comp_v[2][32])
                                        );
                                        
                                        compress_module comp_v_545 (
                                            .x(result[2][33]),
                                            .d(4),
                                            .result(comp_v[2][33])
                                        );
                                        
                                        compress_module comp_v_546 (
                                            .x(result[2][34]),
                                            .d(4),
                                            .result(comp_v[2][34])
                                        );
                                        
                                        compress_module comp_v_547 (
                                            .x(result[2][35]),
                                            .d(4),
                                            .result(comp_v[2][35])
                                        );
                                        
                                        compress_module comp_v_548 (
                                            .x(result[2][36]),
                                            .d(4),
                                            .result(comp_v[2][36])
                                        );
                                        
                                        compress_module comp_v_549 (
                                            .x(result[2][37]),
                                            .d(4),
                                            .result(comp_v[2][37])
                                        );
                                        
                                        compress_module comp_v_550 (
                                            .x(result[2][38]),
                                            .d(4),
                                            .result(comp_v[2][38])
                                        );
                                        
                                        compress_module comp_v_551 (
                                            .x(result[2][39]),
                                            .d(4),
                                            .result(comp_v[2][39])
                                        );
                                        
                                        compress_module comp_v_552 (
                                            .x(result[2][40]),
                                            .d(4),
                                            .result(comp_v[2][40])
                                        );
                                        
                                        compress_module comp_v_553 (
                                            .x(result[2][41]),
                                            .d(4),
                                            .result(comp_v[2][41])
                                        );
                                        
                                        compress_module comp_v_554 (
                                            .x(result[2][42]),
                                            .d(4),
                                            .result(comp_v[2][42])
                                        );
                                        
                                        compress_module comp_v_555 (
                                            .x(result[2][43]),
                                            .d(4),
                                            .result(comp_v[2][43])
                                        );
                                        
                                        compress_module comp_v_556 (
                                            .x(result[2][44]),
                                            .d(4),
                                            .result(comp_v[2][44])
                                        );
                                        
                                        compress_module comp_v_557 (
                                            .x(result[2][45]),
                                            .d(4),
                                            .result(comp_v[2][45])
                                        );
                                        
                                        compress_module comp_v_558 (
                                            .x(result[2][46]),
                                            .d(4),
                                            .result(comp_v[2][46])
                                        );
                                        
                                        compress_module comp_v_559 (
                                            .x(result[2][47]),
                                            .d(4),
                                            .result(comp_v[2][47])
                                        );
                                        
                                        compress_module comp_v_560 (
                                            .x(result[2][48]),
                                            .d(4),
                                            .result(comp_v[2][48])
                                        );
                                        
                                        compress_module comp_v_561 (
                                            .x(result[2][49]),
                                            .d(4),
                                            .result(comp_v[2][49])
                                        );
                                        
                                        compress_module comp_v_562 (
                                            .x(result[2][50]),
                                            .d(4),
                                            .result(comp_v[2][50])
                                        );
                                        
                                        compress_module comp_v_563 (
                                            .x(result[2][51]),
                                            .d(4),
                                            .result(comp_v[2][51])
                                        );
                                        
                                        compress_module comp_v_564 (
                                            .x(result[2][52]),
                                            .d(4),
                                            .result(comp_v[2][52])
                                        );
                                        
                                        compress_module comp_v_565 (
                                            .x(result[2][53]),
                                            .d(4),
                                            .result(comp_v[2][53])
                                        );
                                        
                                        compress_module comp_v_566 (
                                            .x(result[2][54]),
                                            .d(4),
                                            .result(comp_v[2][54])
                                        );
                                        
                                        compress_module comp_v_567 (
                                            .x(result[2][55]),
                                            .d(4),
                                            .result(comp_v[2][55])
                                        );
                                        
                                        compress_module comp_v_568 (
                                            .x(result[2][56]),
                                            .d(4),
                                            .result(comp_v[2][56])
                                        );
                                        
                                        compress_module comp_v_569 (
                                            .x(result[2][57]),
                                            .d(4),
                                            .result(comp_v[2][57])
                                        );
                                        
                                        compress_module comp_v_570 (
                                            .x(result[2][58]),
                                            .d(4),
                                            .result(comp_v[2][58])
                                        );
                                        
                                        compress_module comp_v_571 (
                                            .x(result[2][59]),
                                            .d(4),
                                            .result(comp_v[2][59])
                                        );
                                        
                                        compress_module comp_v_572 (
                                            .x(result[2][60]),
                                            .d(4),
                                            .result(comp_v[2][60])
                                        );
                                        
                                        compress_module comp_v_573 (
                                            .x(result[2][61]),
                                            .d(4),
                                            .result(comp_v[2][61])
                                        );
                                        
                                        compress_module comp_v_574 (
                                            .x(result[2][62]),
                                            .d(4),
                                            .result(comp_v[2][62])
                                        );
                                        
                                        compress_module comp_v_575 (
                                            .x(result[2][63]),
                                            .d(4),
                                            .result(comp_v[2][63])
                                        );
                                        
                                        compress_module comp_v_576 (
                                            .x(result[2][64]),
                                            .d(4),
                                            .result(comp_v[2][64])
                                        );
                                        
                                        compress_module comp_v_577 (
                                            .x(result[2][65]),
                                            .d(4),
                                            .result(comp_v[2][65])
                                        );
                                        
                                        compress_module comp_v_578 (
                                            .x(result[2][66]),
                                            .d(4),
                                            .result(comp_v[2][66])
                                        );
                                        
                                        compress_module comp_v_579 (
                                            .x(result[2][67]),
                                            .d(4),
                                            .result(comp_v[2][67])
                                        );
                                        
                                        compress_module comp_v_580 (
                                            .x(result[2][68]),
                                            .d(4),
                                            .result(comp_v[2][68])
                                        );
                                        
                                        compress_module comp_v_581 (
                                            .x(result[2][69]),
                                            .d(4),
                                            .result(comp_v[2][69])
                                        );
                                        
                                        compress_module comp_v_582 (
                                            .x(result[2][70]),
                                            .d(4),
                                            .result(comp_v[2][70])
                                        );
                                        
                                        compress_module comp_v_583 (
                                            .x(result[2][71]),
                                            .d(4),
                                            .result(comp_v[2][71])
                                        );
                                        
                                        compress_module comp_v_584 (
                                            .x(result[2][72]),
                                            .d(4),
                                            .result(comp_v[2][72])
                                        );
                                        
                                        compress_module comp_v_585 (
                                            .x(result[2][73]),
                                            .d(4),
                                            .result(comp_v[2][73])
                                        );
                                        
                                        compress_module comp_v_586 (
                                            .x(result[2][74]),
                                            .d(4),
                                            .result(comp_v[2][74])
                                        );
                                        
                                        compress_module comp_v_587 (
                                            .x(result[2][75]),
                                            .d(4),
                                            .result(comp_v[2][75])
                                        );
                                        
                                        compress_module comp_v_588 (
                                            .x(result[2][76]),
                                            .d(4),
                                            .result(comp_v[2][76])
                                        );
                                        
                                        compress_module comp_v_589 (
                                            .x(result[2][77]),
                                            .d(4),
                                            .result(comp_v[2][77])
                                        );
                                        
                                        compress_module comp_v_590 (
                                            .x(result[2][78]),
                                            .d(4),
                                            .result(comp_v[2][78])
                                        );
                                        
                                        compress_module comp_v_591 (
                                            .x(result[2][79]),
                                            .d(4),
                                            .result(comp_v[2][79])
                                        );
                                        
                                        compress_module comp_v_592 (
                                            .x(result[2][80]),
                                            .d(4),
                                            .result(comp_v[2][80])
                                        );
                                        
                                        compress_module comp_v_593 (
                                            .x(result[2][81]),
                                            .d(4),
                                            .result(comp_v[2][81])
                                        );
                                        
                                        compress_module comp_v_594 (
                                            .x(result[2][82]),
                                            .d(4),
                                            .result(comp_v[2][82])
                                        );
                                        
                                        compress_module comp_v_595 (
                                            .x(result[2][83]),
                                            .d(4),
                                            .result(comp_v[2][83])
                                        );
                                        
                                        compress_module comp_v_596 (
                                            .x(result[2][84]),
                                            .d(4),
                                            .result(comp_v[2][84])
                                        );
                                        
                                        compress_module comp_v_597 (
                                            .x(result[2][85]),
                                            .d(4),
                                            .result(comp_v[2][85])
                                        );
                                        
                                        compress_module comp_v_598 (
                                            .x(result[2][86]),
                                            .d(4),
                                            .result(comp_v[2][86])
                                        );
                                        
                                        compress_module comp_v_599 (
                                            .x(result[2][87]),
                                            .d(4),
                                            .result(comp_v[2][87])
                                        );
                                        
                                        compress_module comp_v_600 (
                                            .x(result[2][88]),
                                            .d(4),
                                            .result(comp_v[2][88])
                                        );
                                        
                                        compress_module comp_v_601 (
                                            .x(result[2][89]),
                                            .d(4),
                                            .result(comp_v[2][89])
                                        );
                                        
                                        compress_module comp_v_602 (
                                            .x(result[2][90]),
                                            .d(4),
                                            .result(comp_v[2][90])
                                        );
                                        
                                        compress_module comp_v_603 (
                                            .x(result[2][91]),
                                            .d(4),
                                            .result(comp_v[2][91])
                                        );
                                        
                                        compress_module comp_v_604 (
                                            .x(result[2][92]),
                                            .d(4),
                                            .result(comp_v[2][92])
                                        );
                                        
                                        compress_module comp_v_605 (
                                            .x(result[2][93]),
                                            .d(4),
                                            .result(comp_v[2][93])
                                        );
                                        
                                        compress_module comp_v_606 (
                                            .x(result[2][94]),
                                            .d(4),
                                            .result(comp_v[2][94])
                                        );
                                        
                                        compress_module comp_v_607 (
                                            .x(result[2][95]),
                                            .d(4),
                                            .result(comp_v[2][95])
                                        );
                                        
                                        compress_module comp_v_608 (
                                            .x(result[2][96]),
                                            .d(4),
                                            .result(comp_v[2][96])
                                        );
                                        
                                        compress_module comp_v_609 (
                                            .x(result[2][97]),
                                            .d(4),
                                            .result(comp_v[2][97])
                                        );
                                        
                                        compress_module comp_v_610 (
                                            .x(result[2][98]),
                                            .d(4),
                                            .result(comp_v[2][98])
                                        );
                                        
                                        compress_module comp_v_611 (
                                            .x(result[2][99]),
                                            .d(4),
                                            .result(comp_v[2][99])
                                        );
                                        
                                        compress_module comp_v_612 (
                                            .x(result[2][100]),
                                            .d(4),
                                            .result(comp_v[2][100])
                                        );
                                        
                                        compress_module comp_v_613 (
                                            .x(result[2][101]),
                                            .d(4),
                                            .result(comp_v[2][101])
                                        );
                                        
                                        compress_module comp_v_614 (
                                            .x(result[2][102]),
                                            .d(4),
                                            .result(comp_v[2][102])
                                        );
                                        
                                        compress_module comp_v_615 (
                                            .x(result[2][103]),
                                            .d(4),
                                            .result(comp_v[2][103])
                                        );
                                        
                                        compress_module comp_v_616 (
                                            .x(result[2][104]),
                                            .d(4),
                                            .result(comp_v[2][104])
                                        );
                                        
                                        compress_module comp_v_617 (
                                            .x(result[2][105]),
                                            .d(4),
                                            .result(comp_v[2][105])
                                        );
                                        
                                        compress_module comp_v_618 (
                                            .x(result[2][106]),
                                            .d(4),
                                            .result(comp_v[2][106])
                                        );
                                        
                                        compress_module comp_v_619 (
                                            .x(result[2][107]),
                                            .d(4),
                                            .result(comp_v[2][107])
                                        );
                                        
                                        compress_module comp_v_620 (
                                            .x(result[2][108]),
                                            .d(4),
                                            .result(comp_v[2][108])
                                        );
                                        
                                        compress_module comp_v_621 (
                                            .x(result[2][109]),
                                            .d(4),
                                            .result(comp_v[2][109])
                                        );
                                        
                                        compress_module comp_v_622 (
                                            .x(result[2][110]),
                                            .d(4),
                                            .result(comp_v[2][110])
                                        );
                                        
                                        compress_module comp_v_623 (
                                            .x(result[2][111]),
                                            .d(4),
                                            .result(comp_v[2][111])
                                        );
                                        
                                        compress_module comp_v_624 (
                                            .x(result[2][112]),
                                            .d(4),
                                            .result(comp_v[2][112])
                                        );
                                        
                                        compress_module comp_v_625 (
                                            .x(result[2][113]),
                                            .d(4),
                                            .result(comp_v[2][113])
                                        );
                                        
                                        compress_module comp_v_626 (
                                            .x(result[2][114]),
                                            .d(4),
                                            .result(comp_v[2][114])
                                        );
                                        
                                        compress_module comp_v_627 (
                                            .x(result[2][115]),
                                            .d(4),
                                            .result(comp_v[2][115])
                                        );
                                        
                                        compress_module comp_v_628 (
                                            .x(result[2][116]),
                                            .d(4),
                                            .result(comp_v[2][116])
                                        );
                                        
                                        compress_module comp_v_629 (
                                            .x(result[2][117]),
                                            .d(4),
                                            .result(comp_v[2][117])
                                        );
                                        
                                        compress_module comp_v_630 (
                                            .x(result[2][118]),
                                            .d(4),
                                            .result(comp_v[2][118])
                                        );
                                        
                                        compress_module comp_v_631 (
                                            .x(result[2][119]),
                                            .d(4),
                                            .result(comp_v[2][119])
                                        );
                                        
                                        compress_module comp_v_632 (
                                            .x(result[2][120]),
                                            .d(4),
                                            .result(comp_v[2][120])
                                        );
                                        
                                        compress_module comp_v_633 (
                                            .x(result[2][121]),
                                            .d(4),
                                            .result(comp_v[2][121])
                                        );
                                        
                                        compress_module comp_v_634 (
                                            .x(result[2][122]),
                                            .d(4),
                                            .result(comp_v[2][122])
                                        );
                                        
                                        compress_module comp_v_635 (
                                            .x(result[2][123]),
                                            .d(4),
                                            .result(comp_v[2][123])
                                        );
                                        
                                        compress_module comp_v_636 (
                                            .x(result[2][124]),
                                            .d(4),
                                            .result(comp_v[2][124])
                                        );
                                        
                                        compress_module comp_v_637 (
                                            .x(result[2][125]),
                                            .d(4),
                                            .result(comp_v[2][125])
                                        );
                                        
                                        compress_module comp_v_638 (
                                            .x(result[2][126]),
                                            .d(4),
                                            .result(comp_v[2][126])
                                        );
                                        
                                        compress_module comp_v_639 (
                                            .x(result[2][127]),
                                            .d(4),
                                            .result(comp_v[2][127])
                                        );
                                        
                                        compress_module comp_v_640 (
                                            .x(result[2][128]),
                                            .d(4),
                                            .result(comp_v[2][128])
                                        );
                                        
                                        compress_module comp_v_641 (
                                            .x(result[2][129]),
                                            .d(4),
                                            .result(comp_v[2][129])
                                        );
                                        
                                        compress_module comp_v_642 (
                                            .x(result[2][130]),
                                            .d(4),
                                            .result(comp_v[2][130])
                                        );
                                        
                                        compress_module comp_v_643 (
                                            .x(result[2][131]),
                                            .d(4),
                                            .result(comp_v[2][131])
                                        );
                                        
                                        compress_module comp_v_644 (
                                            .x(result[2][132]),
                                            .d(4),
                                            .result(comp_v[2][132])
                                        );
                                        
                                        compress_module comp_v_645 (
                                            .x(result[2][133]),
                                            .d(4),
                                            .result(comp_v[2][133])
                                        );
                                        
                                        compress_module comp_v_646 (
                                            .x(result[2][134]),
                                            .d(4),
                                            .result(comp_v[2][134])
                                        );
                                        
                                        compress_module comp_v_647 (
                                            .x(result[2][135]),
                                            .d(4),
                                            .result(comp_v[2][135])
                                        );
                                        
                                        compress_module comp_v_648 (
                                            .x(result[2][136]),
                                            .d(4),
                                            .result(comp_v[2][136])
                                        );
                                        
                                        compress_module comp_v_649 (
                                            .x(result[2][137]),
                                            .d(4),
                                            .result(comp_v[2][137])
                                        );
                                        
                                        compress_module comp_v_650 (
                                            .x(result[2][138]),
                                            .d(4),
                                            .result(comp_v[2][138])
                                        );
                                        
                                        compress_module comp_v_651 (
                                            .x(result[2][139]),
                                            .d(4),
                                            .result(comp_v[2][139])
                                        );
                                        
                                        compress_module comp_v_652 (
                                            .x(result[2][140]),
                                            .d(4),
                                            .result(comp_v[2][140])
                                        );
                                        
                                        compress_module comp_v_653 (
                                            .x(result[2][141]),
                                            .d(4),
                                            .result(comp_v[2][141])
                                        );
                                        
                                        compress_module comp_v_654 (
                                            .x(result[2][142]),
                                            .d(4),
                                            .result(comp_v[2][142])
                                        );
                                        
                                        compress_module comp_v_655 (
                                            .x(result[2][143]),
                                            .d(4),
                                            .result(comp_v[2][143])
                                        );
                                        
                                        compress_module comp_v_656 (
                                            .x(result[2][144]),
                                            .d(4),
                                            .result(comp_v[2][144])
                                        );
                                        
                                        compress_module comp_v_657 (
                                            .x(result[2][145]),
                                            .d(4),
                                            .result(comp_v[2][145])
                                        );
                                        
                                        compress_module comp_v_658 (
                                            .x(result[2][146]),
                                            .d(4),
                                            .result(comp_v[2][146])
                                        );
                                        
                                        compress_module comp_v_659 (
                                            .x(result[2][147]),
                                            .d(4),
                                            .result(comp_v[2][147])
                                        );
                                        
                                        compress_module comp_v_660 (
                                            .x(result[2][148]),
                                            .d(4),
                                            .result(comp_v[2][148])
                                        );
                                        
                                        compress_module comp_v_661 (
                                            .x(result[2][149]),
                                            .d(4),
                                            .result(comp_v[2][149])
                                        );
                                        
                                        compress_module comp_v_662 (
                                            .x(result[2][150]),
                                            .d(4),
                                            .result(comp_v[2][150])
                                        );
                                        
                                        compress_module comp_v_663 (
                                            .x(result[2][151]),
                                            .d(4),
                                            .result(comp_v[2][151])
                                        );
                                        
                                        compress_module comp_v_664 (
                                            .x(result[2][152]),
                                            .d(4),
                                            .result(comp_v[2][152])
                                        );
                                        
                                        compress_module comp_v_665 (
                                            .x(result[2][153]),
                                            .d(4),
                                            .result(comp_v[2][153])
                                        );
                                        
                                        compress_module comp_v_666 (
                                            .x(result[2][154]),
                                            .d(4),
                                            .result(comp_v[2][154])
                                        );
                                        
                                        compress_module comp_v_667 (
                                            .x(result[2][155]),
                                            .d(4),
                                            .result(comp_v[2][155])
                                        );
                                        
                                        compress_module comp_v_668 (
                                            .x(result[2][156]),
                                            .d(4),
                                            .result(comp_v[2][156])
                                        );
                                        
                                        compress_module comp_v_669 (
                                            .x(result[2][157]),
                                            .d(4),
                                            .result(comp_v[2][157])
                                        );
                                        
                                        compress_module comp_v_670 (
                                            .x(result[2][158]),
                                            .d(4),
                                            .result(comp_v[2][158])
                                        );
                                        
                                        compress_module comp_v_671 (
                                            .x(result[2][159]),
                                            .d(4),
                                            .result(comp_v[2][159])
                                        );
                                        
                                        compress_module comp_v_672 (
                                            .x(result[2][160]),
                                            .d(4),
                                            .result(comp_v[2][160])
                                        );
                                        
                                        compress_module comp_v_673 (
                                            .x(result[2][161]),
                                            .d(4),
                                            .result(comp_v[2][161])
                                        );
                                        
                                        compress_module comp_v_674 (
                                            .x(result[2][162]),
                                            .d(4),
                                            .result(comp_v[2][162])
                                        );
                                        
                                        compress_module comp_v_675 (
                                            .x(result[2][163]),
                                            .d(4),
                                            .result(comp_v[2][163])
                                        );
                                        
                                        compress_module comp_v_676 (
                                            .x(result[2][164]),
                                            .d(4),
                                            .result(comp_v[2][164])
                                        );
                                        
                                        compress_module comp_v_677 (
                                            .x(result[2][165]),
                                            .d(4),
                                            .result(comp_v[2][165])
                                        );
                                        
                                        compress_module comp_v_678 (
                                            .x(result[2][166]),
                                            .d(4),
                                            .result(comp_v[2][166])
                                        );
                                        
                                        compress_module comp_v_679 (
                                            .x(result[2][167]),
                                            .d(4),
                                            .result(comp_v[2][167])
                                        );
                                        
                                        compress_module comp_v_680 (
                                            .x(result[2][168]),
                                            .d(4),
                                            .result(comp_v[2][168])
                                        );
                                        
                                        compress_module comp_v_681 (
                                            .x(result[2][169]),
                                            .d(4),
                                            .result(comp_v[2][169])
                                        );
                                        
                                        compress_module comp_v_682 (
                                            .x(result[2][170]),
                                            .d(4),
                                            .result(comp_v[2][170])
                                        );
                                        
                                        compress_module comp_v_683 (
                                            .x(result[2][171]),
                                            .d(4),
                                            .result(comp_v[2][171])
                                        );
                                        
                                        compress_module comp_v_684 (
                                            .x(result[2][172]),
                                            .d(4),
                                            .result(comp_v[2][172])
                                        );
                                        
                                        compress_module comp_v_685 (
                                            .x(result[2][173]),
                                            .d(4),
                                            .result(comp_v[2][173])
                                        );
                                        
                                        compress_module comp_v_686 (
                                            .x(result[2][174]),
                                            .d(4),
                                            .result(comp_v[2][174])
                                        );
                                        
                                        compress_module comp_v_687 (
                                            .x(result[2][175]),
                                            .d(4),
                                            .result(comp_v[2][175])
                                        );
                                        
                                        compress_module comp_v_688 (
                                            .x(result[2][176]),
                                            .d(4),
                                            .result(comp_v[2][176])
                                        );
                                        
                                        compress_module comp_v_689 (
                                            .x(result[2][177]),
                                            .d(4),
                                            .result(comp_v[2][177])
                                        );
                                        
                                        compress_module comp_v_690 (
                                            .x(result[2][178]),
                                            .d(4),
                                            .result(comp_v[2][178])
                                        );
                                        
                                        compress_module comp_v_691 (
                                            .x(result[2][179]),
                                            .d(4),
                                            .result(comp_v[2][179])
                                        );
                                        
                                        compress_module comp_v_692 (
                                            .x(result[2][180]),
                                            .d(4),
                                            .result(comp_v[2][180])
                                        );
                                        
                                        compress_module comp_v_693 (
                                            .x(result[2][181]),
                                            .d(4),
                                            .result(comp_v[2][181])
                                        );
                                        
                                        compress_module comp_v_694 (
                                            .x(result[2][182]),
                                            .d(4),
                                            .result(comp_v[2][182])
                                        );
                                        
                                        compress_module comp_v_695 (
                                            .x(result[2][183]),
                                            .d(4),
                                            .result(comp_v[2][183])
                                        );
                                        
                                        compress_module comp_v_696 (
                                            .x(result[2][184]),
                                            .d(4),
                                            .result(comp_v[2][184])
                                        );
                                        
                                        compress_module comp_v_697 (
                                            .x(result[2][185]),
                                            .d(4),
                                            .result(comp_v[2][185])
                                        );
                                        
                                        compress_module comp_v_698 (
                                            .x(result[2][186]),
                                            .d(4),
                                            .result(comp_v[2][186])
                                        );
                                        
                                        compress_module comp_v_699 (
                                            .x(result[2][187]),
                                            .d(4),
                                            .result(comp_v[2][187])
                                        );
                                        
                                        compress_module comp_v_700 (
                                            .x(result[2][188]),
                                            .d(4),
                                            .result(comp_v[2][188])
                                        );
                                        
                                        compress_module comp_v_701 (
                                            .x(result[2][189]),
                                            .d(4),
                                            .result(comp_v[2][189])
                                        );
                                        
                                        compress_module comp_v_702 (
                                            .x(result[2][190]),
                                            .d(4),
                                            .result(comp_v[2][190])
                                        );
                                        
                                        compress_module comp_v_703 (
                                            .x(result[2][191]),
                                            .d(4),
                                            .result(comp_v[2][191])
                                        );
                                        
                                        compress_module comp_v_704 (
                                            .x(result[2][192]),
                                            .d(4),
                                            .result(comp_v[2][192])
                                        );
                                        
                                        compress_module comp_v_705 (
                                            .x(result[2][193]),
                                            .d(4),
                                            .result(comp_v[2][193])
                                        );
                                        
                                        compress_module comp_v_706 (
                                            .x(result[2][194]),
                                            .d(4),
                                            .result(comp_v[2][194])
                                        );
                                        
                                        compress_module comp_v_707 (
                                            .x(result[2][195]),
                                            .d(4),
                                            .result(comp_v[2][195])
                                        );
                                        
                                        compress_module comp_v_708 (
                                            .x(result[2][196]),
                                            .d(4),
                                            .result(comp_v[2][196])
                                        );
                                        
                                        compress_module comp_v_709 (
                                            .x(result[2][197]),
                                            .d(4),
                                            .result(comp_v[2][197])
                                        );
                                        
                                        compress_module comp_v_710 (
                                            .x(result[2][198]),
                                            .d(4),
                                            .result(comp_v[2][198])
                                        );
                                        
                                        compress_module comp_v_711 (
                                            .x(result[2][199]),
                                            .d(4),
                                            .result(comp_v[2][199])
                                        );
                                        
                                        compress_module comp_v_712 (
                                            .x(result[2][200]),
                                            .d(4),
                                            .result(comp_v[2][200])
                                        );
                                        
                                        compress_module comp_v_713 (
                                            .x(result[2][201]),
                                            .d(4),
                                            .result(comp_v[2][201])
                                        );
                                        
                                        compress_module comp_v_714 (
                                            .x(result[2][202]),
                                            .d(4),
                                            .result(comp_v[2][202])
                                        );
                                        
                                        compress_module comp_v_715 (
                                            .x(result[2][203]),
                                            .d(4),
                                            .result(comp_v[2][203])
                                        );
                                        
                                        compress_module comp_v_716 (
                                            .x(result[2][204]),
                                            .d(4),
                                            .result(comp_v[2][204])
                                        );
                                        
                                        compress_module comp_v_717 (
                                            .x(result[2][205]),
                                            .d(4),
                                            .result(comp_v[2][205])
                                        );
                                        
                                        compress_module comp_v_718 (
                                            .x(result[2][206]),
                                            .d(4),
                                            .result(comp_v[2][206])
                                        );
                                        
                                        compress_module comp_v_719 (
                                            .x(result[2][207]),
                                            .d(4),
                                            .result(comp_v[2][207])
                                        );
                                        
                                        compress_module comp_v_720 (
                                            .x(result[2][208]),
                                            .d(4),
                                            .result(comp_v[2][208])
                                        );
                                        
                                        compress_module comp_v_721 (
                                            .x(result[2][209]),
                                            .d(4),
                                            .result(comp_v[2][209])
                                        );
                                        
                                        compress_module comp_v_722 (
                                            .x(result[2][210]),
                                            .d(4),
                                            .result(comp_v[2][210])
                                        );
                                        
                                        compress_module comp_v_723 (
                                            .x(result[2][211]),
                                            .d(4),
                                            .result(comp_v[2][211])
                                        );
                                        
                                        compress_module comp_v_724 (
                                            .x(result[2][212]),
                                            .d(4),
                                            .result(comp_v[2][212])
                                        );
                                        
                                        compress_module comp_v_725 (
                                            .x(result[2][213]),
                                            .d(4),
                                            .result(comp_v[2][213])
                                        );
                                        
                                        compress_module comp_v_726 (
                                            .x(result[2][214]),
                                            .d(4),
                                            .result(comp_v[2][214])
                                        );
                                        
                                        compress_module comp_v_727 (
                                            .x(result[2][215]),
                                            .d(4),
                                            .result(comp_v[2][215])
                                        );
                                        
                                        compress_module comp_v_728 (
                                            .x(result[2][216]),
                                            .d(4),
                                            .result(comp_v[2][216])
                                        );
                                        
                                        compress_module comp_v_729 (
                                            .x(result[2][217]),
                                            .d(4),
                                            .result(comp_v[2][217])
                                        );
                                        
                                        compress_module comp_v_730 (
                                            .x(result[2][218]),
                                            .d(4),
                                            .result(comp_v[2][218])
                                        );
                                        
                                        compress_module comp_v_731 (
                                            .x(result[2][219]),
                                            .d(4),
                                            .result(comp_v[2][219])
                                        );
                                        
                                        compress_module comp_v_732 (
                                            .x(result[2][220]),
                                            .d(4),
                                            .result(comp_v[2][220])
                                        );
                                        
                                        compress_module comp_v_733 (
                                            .x(result[2][221]),
                                            .d(4),
                                            .result(comp_v[2][221])
                                        );
                                        
                                        compress_module comp_v_734 (
                                            .x(result[2][222]),
                                            .d(4),
                                            .result(comp_v[2][222])
                                        );
                                        
                                        compress_module comp_v_735 (
                                            .x(result[2][223]),
                                            .d(4),
                                            .result(comp_v[2][223])
                                        );
                                        
                                        compress_module comp_v_736 (
                                            .x(result[2][224]),
                                            .d(4),
                                            .result(comp_v[2][224])
                                        );
                                        
                                        compress_module comp_v_737 (
                                            .x(result[2][225]),
                                            .d(4),
                                            .result(comp_v[2][225])
                                        );
                                        
                                        compress_module comp_v_738 (
                                            .x(result[2][226]),
                                            .d(4),
                                            .result(comp_v[2][226])
                                        );
                                        
                                        compress_module comp_v_739 (
                                            .x(result[2][227]),
                                            .d(4),
                                            .result(comp_v[2][227])
                                        );
                                        
                                        compress_module comp_v_740 (
                                            .x(result[2][228]),
                                            .d(4),
                                            .result(comp_v[2][228])
                                        );
                                        
                                        compress_module comp_v_741 (
                                            .x(result[2][229]),
                                            .d(4),
                                            .result(comp_v[2][229])
                                        );
                                        
                                        compress_module comp_v_742 (
                                            .x(result[2][230]),
                                            .d(4),
                                            .result(comp_v[2][230])
                                        );
                                        
                                        compress_module comp_v_743 (
                                            .x(result[2][231]),
                                            .d(4),
                                            .result(comp_v[2][231])
                                        );
                                        
                                        compress_module comp_v_744 (
                                            .x(result[2][232]),
                                            .d(4),
                                            .result(comp_v[2][232])
                                        );
                                        
                                        compress_module comp_v_745 (
                                            .x(result[2][233]),
                                            .d(4),
                                            .result(comp_v[2][233])
                                        );
                                        
                                        compress_module comp_v_746 (
                                            .x(result[2][234]),
                                            .d(4),
                                            .result(comp_v[2][234])
                                        );
                                        
                                        compress_module comp_v_747 (
                                            .x(result[2][235]),
                                            .d(4),
                                            .result(comp_v[2][235])
                                        );
                                        
                                        compress_module comp_v_748 (
                                            .x(result[2][236]),
                                            .d(4),
                                            .result(comp_v[2][236])
                                        );
                                        
                                        compress_module comp_v_749 (
                                            .x(result[2][237]),
                                            .d(4),
                                            .result(comp_v[2][237])
                                        );
                                        
                                        compress_module comp_v_750 (
                                            .x(result[2][238]),
                                            .d(4),
                                            .result(comp_v[2][238])
                                        );
                                        
                                        compress_module comp_v_751 (
                                            .x(result[2][239]),
                                            .d(4),
                                            .result(comp_v[2][239])
                                        );
                                        
                                        compress_module comp_v_752 (
                                            .x(result[2][240]),
                                            .d(4),
                                            .result(comp_v[2][240])
                                        );
                                        
                                        compress_module comp_v_753 (
                                            .x(result[2][241]),
                                            .d(4),
                                            .result(comp_v[2][241])
                                        );
                                        
                                        compress_module comp_v_754 (
                                            .x(result[2][242]),
                                            .d(4),
                                            .result(comp_v[2][242])
                                        );
                                        
                                        compress_module comp_v_755 (
                                            .x(result[2][243]),
                                            .d(4),
                                            .result(comp_v[2][243])
                                        );
                                        
                                        compress_module comp_v_756 (
                                            .x(result[2][244]),
                                            .d(4),
                                            .result(comp_v[2][244])
                                        );
                                        
                                        compress_module comp_v_757 (
                                            .x(result[2][245]),
                                            .d(4),
                                            .result(comp_v[2][245])
                                        );
                                        
                                        compress_module comp_v_758 (
                                            .x(result[2][246]),
                                            .d(4),
                                            .result(comp_v[2][246])
                                        );
                                        
                                        compress_module comp_v_759 (
                                            .x(result[2][247]),
                                            .d(4),
                                            .result(comp_v[2][247])
                                        );
                                        
                                        compress_module comp_v_760 (
                                            .x(result[2][248]),
                                            .d(4),
                                            .result(comp_v[2][248])
                                        );
                                        
                                        compress_module comp_v_761 (
                                            .x(result[2][249]),
                                            .d(4),
                                            .result(comp_v[2][249])
                                        );
                                        
                                        compress_module comp_v_762 (
                                            .x(result[2][250]),
                                            .d(4),
                                            .result(comp_v[2][250])
                                        );
                                        
                                        compress_module comp_v_763 (
                                            .x(result[2][251]),
                                            .d(4),
                                            .result(comp_v[2][251])
                                        );
                                        
                                        compress_module comp_v_764 (
                                            .x(result[2][252]),
                                            .d(4),
                                            .result(comp_v[2][252])
                                        );
                                        
                                        compress_module comp_v_765 (
                                            .x(result[2][253]),
                                            .d(4),
                                            .result(comp_v[2][253])
                                        );
                                        
                                        compress_module comp_v_766 (
                                            .x(result[2][254]),
                                            .d(4),
                                            .result(comp_v[2][254])
                                        );
                                        
                                        compress_module comp_v_767 (
                                            .x(result[2][255]),
                                            .d(4),
                                            .result(comp_v[2][255])
                                        );
                                          
                                        encode #(.D(8),.BYTE_LEN(32))enc_u0 (
                                            .F(com_out[0]),
                                            .B(encode_u[0])
                                        );
                                        
                                        encode #(.D(8),.BYTE_LEN(32))enc_u1 (
                                            .F(com_out[1]),
                                            .B(encode_u[1])
                                        );
                                        
                                        encode #(.D(8),.BYTE_LEN(32))enc_u2 (
                                            .F(com_out[2]),
                                            .B(encode_u[2])
                                        );
                                        encode #(.D(8),.BYTE_LEN(32))enc_v0 (
                                            .F(comp_v[0]),
                                            .B(encode_v[0])
                                        );
                                        
                                        encode #(.D(8),.BYTE_LEN(32))enc_v1 (
                                            .F(comp_v[1]),
                                            .B(encode_v[1])
                                        );
                                        
                                        encode #(.D(8),.BYTE_LEN(32))enc_v2 (
                                            .F(comp_v[2]),
                                            .B(encode_v[2])
                                        );
                                        
always_ff @(posedge clk or posedge rst) begin
                                     if (rst) begin
                                     ntt_started <=0;
                                         all_shake_done <= 0;
                                         mul <= 0;
                          //                       start_encode <= 0;
                                                 start_parse  <= 0;
                                                 start_cbd    <= 0;
                                                 start_prf    <= 0;
                          //                       start_ntt <= 0;
                                     end else begin
                          //           start_mul <=0;
                          //           start_encode<=0;
                          //ntt_started <=0;
//                          start_ntt <= 0;
                          
//                                     start_mul    <= 0;
                          //                   start_encode <= 0;
                                             start_parse  <= 0;
                                             start_cbd    <= 0;
                                             start_prf    <= 0;
                                      start1 <= 1;
                                     zetas[0] = 17; zetas[1] = 2761; zetas[2] = 583; zetas[3] = 2649; zetas[4] = 1637; zetas[5] = 723; zetas[6] = 2288; zetas[7] = 1100;
                                             zetas[8] = 1409; zetas[9] = 2662; zetas[10] = 3281; zetas[11] = 233; zetas[12] = 756; zetas[13] = 2156; zetas[14] = 3015; zetas[15] = 3050;
                                             zetas[16] = 1703; zetas[17] = 1651; zetas[18] = 2789; zetas[19] = 1789; zetas[20] = 1847; zetas[21] = 952; zetas[22] = 1461; zetas[23] = 2687;
                                             zetas[24] = 939; zetas[25] = 2308; zetas[26] = 2437; zetas[27] = 2388; zetas[28] = 733; zetas[29] = 2337; zetas[30] = 268; zetas[31] = 641;
                                             zetas[32] = 1584; zetas[33] = 2298; zetas[34] = 2037; zetas[35] = 3220; zetas[36] = 375; zetas[37] = 2549; zetas[38] = 2090; zetas[39] = 1645;
                                             zetas[40] = 1063; zetas[41] = 319; zetas[42] = 2773; zetas[43] = 757; zetas[44] = 2099; zetas[45] = 561; zetas[46] = 2466; zetas[47] = 2594;
                                             zetas[48] = 2804; zetas[49] = 1092; zetas[50] = 403; zetas[51] = 1026; zetas[52] = 1143; zetas[53] = 2150; zetas[54] = 2775; zetas[55] = 886;
                                             zetas[56] = 1722; zetas[57] = 1212; zetas[58] = 1874; zetas[59] = 1029; zetas[60] = 2110; zetas[61] = 2935; zetas[62] = 885; zetas[63] = 2154;
                                             zetas[64] = 289; zetas[65] = 331; zetas[66] = 3253; zetas[67] = 1756; zetas[68] = 1197; zetas[69] = 2304; zetas[70] = 2277; zetas[71] = 2055;
                                             zetas[72] = 650; zetas[73] = 1977; zetas[74] = 2513; zetas[75] = 632; zetas[76] = 2865; zetas[77] = 33; zetas[78] = 1320; zetas[79] = 1915;
                                             zetas[80] = 2319; zetas[81] = 1435; zetas[82] = 807; zetas[83] = 452; zetas[84] = 1438; zetas[85] = 2868; zetas[86] = 1534; zetas[87] = 2402;
                                             zetas[88] = 2647; zetas[89] = 2617; zetas[90] = 1481; zetas[91] = 648; zetas[92] = 2474; zetas[93] = 3110; zetas[94] = 1227; zetas[95] = 910;
                                             zetas[96] = 296; zetas[97] = 2447; zetas[98] = 1339; zetas[99] = 1476; zetas[100] = 3046; zetas[101] = 56; zetas[102] = 2240; zetas[103] = 1333;
                                             zetas[104] = 1426; zetas[105] = 2094; zetas[106] = 535; zetas[107] = 2882; zetas[108] = 2393; zetas[109] = 2879; zetas[110] = 1974; zetas[111] = 821;
                                             zetas[112] = 1062; zetas[113] = 1919; zetas[114] = 193; zetas[115] = 797; zetas[116] = 2786; zetas[117] = 3260; zetas[118] = 569; zetas[119] = 1746;
                                             zetas[120] = 2642; zetas[121] = 630; zetas[122] = 1897; zetas[123] = 848; zetas[124] = 2580; zetas[125] = 3289; zetas[126] = 1729; zetas[127] = 3328;
                                      zetas[17] = 2637;
                                   
                                   
                                    for (int i = 0; i < 768; i = i + 1) begin
                                                     
                                                                    parse_array1[i] = xof[(i+1)*8-1 -: 8];
                                                                     parse_array2[i] = xof2[(i+1)*8-1 -: 8];
                                                                      parse_array3[i] = xof3[(i+1)*8-1 -: 8];
                                                                       parse_array4[i] = xof4[(i+1)*8-1 -: 8];
                                                                        parse_array5[i] = xof5[(i+1)*8-1 -: 8];
                                                                         parse_array6[i] = xof6[(i+1)*8-1 -: 8];
                                                                          parse_array7[i] = xof7[(i+1)*8-1 -: 8];
                                                                           parse_array8[i] = xof8[(i+1)*8-1 -: 8];
                                                                            parse_array9[i] = xof9[(i+1)*8-1 -: 8];
                                                                       
                                     end
                                      if (done0_shake && done1_shake && done2_shake && done3_shake
                                                       && done6_shake && done7_shake && done8_shake  ) begin
                                                       start_parse <= 1;
                                                       start1 <= 0; 
                                                   end
                                                   
                                      if (done0 && done1 && done2 && done3 && done4 && done5 && done6 && done7 && done8 && !done9_shake && !done10_shake && !done11_shake && !done12_shake && !done13_shake && !done14_shake) begin
                                                                                start_parse <= 0;
                                                                                start_prf <= 1;
                                                                                 
                                                                            end
                            for (int i = 0; i < 128; i++) begin
                                                       prf_bytes_0[i] = prf_0[8*i +: 8];
                                                       prf_bytes_1[i] = prf_1[8*i +: 8];
                                                       prf_bytes_2[i] = prf_2[8*i +: 8];
                                                       prf_bytes_3[i] = prf_3[8*i +: 8];
                                                       prf_bytes_4[i] = prf_4[8*i +: 8];
                                                       prf_bytes_5[i] = prf_5[8*i +: 8];
                                                       prf_bytes_6[i] = prf_6[8*i +: 8];
                                                   end
                          //            
                                            if (done0_shake && done1_shake && done2_shake && done3_shake &&
                                                done4_shake && done5_shake && done6_shake && done7_shake && done8_shake) begin
                                                all_shake_done <= 1;
                                                start1 <= 0; 
                                            end else begin
                                                all_shake_done <= 0; 
                                            end
                                       
                                             if (done0_mul && done1_mul && done2_mul && done3_mul && done4_mul && done5_mul && done6_mul && done7_mul && done8_mul) begin
                                                                                                                                           mul_add[0][0] <= ((mult_out_00[0] + mult_out_01[0] + mult_out_02[0])%3329);
                                                                                                                                           mul_add[0][1] <= ((mult_out_00[1] + mult_out_01[1] + mult_out_02[1])%3329) ;
                                                                                                                                           mul_add[0][2] <= ((mult_out_00[2] + mult_out_01[2] + mult_out_02[2])%3329) ;
                                                                                                                                           mul_add[0][3] <= ((mult_out_00[3] + mult_out_01[3] + mult_out_02[3])%3329) ;
                                                                                                                                           mul_add[0][4] <= ((mult_out_00[4] + mult_out_01[4] + mult_out_02[4])%3329) ;
                                                                                                                                           mul_add[0][5]<=((mult_out_00[5] + mult_out_01[5] + mult_out_02[5])%3329) ;
                                                                                                                                           mul_add[0][6]<=((mult_out_00[6] + mult_out_01[6] + mult_out_02[6])%3329);
                                                                                                                                           mul_add[0][7]<=((mult_out_00[7] + mult_out_01[7] + mult_out_02[7])%3329) ;
                                                                                                                                           mul_add[0][8]<=((mult_out_00[8] + mult_out_01[8] + mult_out_02[8])%3329);
                                                                                                                                           mul_add[0][9]<=((mult_out_00[9] + mult_out_01[9] + mult_out_02[9])%3329) ;
                                                                                                                                           mul_add[0][10]<=((mult_out_00[10] + mult_out_01[10] + mult_out_02[10])%3329) ;
                                                                                                                                           mul_add[0][11]<=((mult_out_00[11] + mult_out_01[11] + mult_out_02[11])%3329) ;
                                                                                                                                           mul_add[0][12]<=((mult_out_00[12] + mult_out_01[12] + mult_out_02[12])%3329) ;
                                                                                                                                           mul_add[0][13]<=((mult_out_00[13] + mult_out_01[13] + mult_out_02[13])%3329) ;
                                                                                                                                           mul_add[0][14]<=((mult_out_00[14] + mult_out_01[14] + mult_out_02[14])%3329) ;
                                                                                                                                           mul_add[0][15]<=((mult_out_00[15] + mult_out_01[15] + mult_out_02[15])%3329) ;
                                                                                                                                           mul_add[0][16]<=((mult_out_00[16] + mult_out_01[16] + mult_out_02[16])%3329) ;
                                                                                                                                           mul_add[0][17]<=((mult_out_00[17] + mult_out_01[17] + mult_out_02[17])%3329) ;
                                                                                                                                           mul_add[0][18]<=((mult_out_00[18] + mult_out_01[18] + mult_out_02[18])%3329) ;
                                                                                                                                           mul_add[0][19]<=((mult_out_00[19] + mult_out_01[19] + mult_out_02[19])%3329) ;
                                                                                                                                           mul_add[0][20]<=((mult_out_00[20] + mult_out_01[20] + mult_out_02[20])%3329) ;
                                                                                                                                           mul_add[0][21]<=((mult_out_00[21] + mult_out_01[21] + mult_out_02[21])%3329) ;
                                                                                                                                           mul_add[0][22]<=((mult_out_00[22] + mult_out_01[22] + mult_out_02[22])%3329) ;
                                                                                                                                           mul_add[0][23]<=((mult_out_00[23] + mult_out_01[23] + mult_out_02[23])%3329) ;
                                                                                                                                           mul_add[0][24]<=((mult_out_00[24] + mult_out_01[24] + mult_out_02[24])%3329) ;
                                                                                                                                           mul_add[0][25]<=((mult_out_00[25] + mult_out_01[25] + mult_out_02[25])%3329) ;
                                                                                                                                           mul_add[0][26]<=((mult_out_00[26] + mult_out_01[26] + mult_out_02[26])%3329) ;
                                                                                                                                           mul_add[0][27]<=((mult_out_00[27] + mult_out_01[27] + mult_out_02[27])%3329) ;
                                                                                                                                           mul_add[0][28]<=((mult_out_00[28] + mult_out_01[28] + mult_out_02[28])%3329) ;
                                                                                                                                           mul_add[0][29]<=((mult_out_00[29] + mult_out_01[29] + mult_out_02[29])%3329) ;
                                                                                                                                           mul_add[0][30]<=((mult_out_00[30] + mult_out_01[30] + mult_out_02[30])%3329) ;
                                                                                                                                           mul_add[0][31]<=((mult_out_00[31] + mult_out_01[31] + mult_out_02[31])%3329) ;
                                                                                                                                           mul_add[0][32]<=((mult_out_00[32] + mult_out_01[32] + mult_out_02[32])%3329) ;
                                                                                                                                           mul_add[0][33]<=((mult_out_00[33] + mult_out_01[33] + mult_out_02[33])%3329) ;
                                                                                                                                           mul_add[0][34]<=((mult_out_00[34] + mult_out_01[34] + mult_out_02[34])%3329) ;
                                                                                                                                           mul_add[0][35]<=((mult_out_00[35] + mult_out_01[35] + mult_out_02[35])%3329) ;
                                                                                                                                           mul_add[0][36]<=((mult_out_00[36] + mult_out_01[36] + mult_out_02[36])%3329) ;
                                                                                                                                           mul_add[0][37]<=((mult_out_00[37] + mult_out_01[37] + mult_out_02[37])%3329) ;
                                                                                                                                           mul_add[0][38]<=((mult_out_00[38] + mult_out_01[38] + mult_out_02[38])%3329) ;
                                                                                                                                           mul_add[0][39]<=((mult_out_00[39] + mult_out_01[39] + mult_out_02[39])%3329) ;
                                                                                                                                           mul_add[0][40]<=((mult_out_00[40] + mult_out_01[40] + mult_out_02[40])%3329) ;
                                                                                                                                           mul_add[0][41]<=((mult_out_00[41] + mult_out_01[41] + mult_out_02[41])%3329) ;
                                                                                                                                           mul_add[0][42]<=((mult_out_00[42] + mult_out_01[42] + mult_out_02[42])%3329) ;
                                                                                                                                           mul_add[0][43]<=((mult_out_00[43] + mult_out_01[43] + mult_out_02[43])%3329) ;
                                                                                                                                           mul_add[0][44]<=((mult_out_00[44] + mult_out_01[44] + mult_out_02[44])%3329) ;
                                                                                                                                           mul_add[0][45]<=((mult_out_00[45] + mult_out_01[45] + mult_out_02[45])%3329) ;
                                                                                                                                           mul_add[0][46]<=((mult_out_00[46] + mult_out_01[46] + mult_out_02[46])%3329) ;
                                                                                                                                           mul_add[0][47]<=((mult_out_00[47] + mult_out_01[47] + mult_out_02[47])%3329) ;
                                                                                                                                           mul_add[0][48]<=((mult_out_00[48] + mult_out_01[48] + mult_out_02[48])%3329) ;
                                                                                                                                           mul_add[0][49]<=((mult_out_00[49] + mult_out_01[49] + mult_out_02[49])%3329) ;
                                                                                                                                           mul_add[0][50]<=((mult_out_00[50] + mult_out_01[50] + mult_out_02[50])%3329) ;
                                                                                                                                           mul_add[0][51]<=((mult_out_00[51] + mult_out_01[51] + mult_out_02[51])%3329) ;
                                                                                                                                           mul_add[0][52]<=((mult_out_00[52] + mult_out_01[52] + mult_out_02[52])%3329) ;
                                                                                                                                           mul_add[0][53]<=((mult_out_00[53] + mult_out_01[53] + mult_out_02[53])%3329) ;
                                                                                                                                           mul_add[0][54]<=((mult_out_00[54] + mult_out_01[54] + mult_out_02[54])%3329) ;
                                                                                                                                           mul_add[0][55]<=((mult_out_00[55] + mult_out_01[55] + mult_out_02[55])%3329) ;
                                                                                                                                           mul_add[0][56]<=((mult_out_00[56] + mult_out_01[56] + mult_out_02[56])%3329) ;
                                                                                                                                           mul_add[0][57]<=((mult_out_00[57] + mult_out_01[57] + mult_out_02[57])%3329) ;
                                                                                                                                           mul_add[0][58]<=((mult_out_00[58] + mult_out_01[58] + mult_out_02[58])%3329) ;
                                                                                                                                           mul_add[0][59]<=((mult_out_00[59] + mult_out_01[59] + mult_out_02[59])%3329) ;
                                                                                                                                           mul_add[0][60]<=((mult_out_00[60] + mult_out_01[60] + mult_out_02[60])%3329) ;
                                                                                                                                           mul_add[0][61]<=((mult_out_00[61] + mult_out_01[61] + mult_out_02[61])%3329) ;
                                                                                                                                           mul_add[0][62]<=((mult_out_00[62] + mult_out_01[62] + mult_out_02[62])%3329) ;
                                                                                                                                           mul_add[0][63]<=((mult_out_00[63] + mult_out_01[63] + mult_out_02[63])%3329) ;
                                                                                                                                           mul_add[0][64]<=((mult_out_00[64] + mult_out_01[64] + mult_out_02[64])%3329) ;
                                                                                                                                           mul_add[0][65]<=((mult_out_00[65] + mult_out_01[65] + mult_out_02[65])%3329) ;
                                                                                                                                           mul_add[0][66]<=((mult_out_00[66] + mult_out_01[66] + mult_out_02[66])%3329) ;
                                                                                                                                           mul_add[0][67]<=((mult_out_00[67] + mult_out_01[67] + mult_out_02[67])%3329) ;
                                                                                                                                           mul_add[0][68]<=((mult_out_00[68] + mult_out_01[68] + mult_out_02[68])%3329) ;
                                                                                                                                           mul_add[0][69]<=((mult_out_00[69] + mult_out_01[69] + mult_out_02[69])%3329) ;
                                                                                                                                           mul_add[0][70]<=((mult_out_00[70] + mult_out_01[70] + mult_out_02[70])%3329) ;
                                                                                                                                           mul_add[0][71]<=((mult_out_00[71] + mult_out_01[71] + mult_out_02[71])%3329) ;
                                                                                                                                           mul_add[0][72]<=((mult_out_00[72] + mult_out_01[72] + mult_out_02[72])%3329) ;
                                                                                                                                           mul_add[0][73]<=((mult_out_00[73] + mult_out_01[73] + mult_out_02[73])%3329) ;
                                                                                                                                           mul_add[0][74]<=((mult_out_00[74] + mult_out_01[74] + mult_out_02[74])%3329) ;
                                                                                                                                           mul_add[0][75]<=((mult_out_00[75] + mult_out_01[75] + mult_out_02[75])%3329) ;
                                                                                                                                           mul_add[0][76]<=((mult_out_00[76] + mult_out_01[76] + mult_out_02[76])%3329) ;
                                                                                                                                           mul_add[0][77]<=((mult_out_00[77] + mult_out_01[77] + mult_out_02[77])%3329) ;
                                                                                                                                           mul_add[0][78]<=((mult_out_00[78] + mult_out_01[78] + mult_out_02[78])%3329) ;
                                                                                                                                           mul_add[0][79]<=((mult_out_00[79] + mult_out_01[79] + mult_out_02[79])%3329) ;
                                                                                                                                           mul_add[0][80]<=((mult_out_00[80] + mult_out_01[80] + mult_out_02[80])%3329) ;
                                                                                                                                           mul_add[0][81]<=((mult_out_00[81] + mult_out_01[81] + mult_out_02[81])%3329) ;
                                                                                                                                           mul_add[0][82]<=((mult_out_00[82] + mult_out_01[82] + mult_out_02[82])%3329) ;
                                                                                                                                           mul_add[0][83]<=((mult_out_00[83] + mult_out_01[83] + mult_out_02[83])%3329) ;
                                                                                                                                           mul_add[0][84]<=((mult_out_00[84] + mult_out_01[84] + mult_out_02[84])%3329) ;
                                                                                                                                           mul_add[0][85]<=((mult_out_00[85] + mult_out_01[85] + mult_out_02[85])%3329) ;
                                                                                                                                           mul_add[0][86]<=((mult_out_00[86] + mult_out_01[86] + mult_out_02[86])%3329) ;
                                                                                                                                           mul_add[0][87]<=((mult_out_00[87] + mult_out_01[87] + mult_out_02[87])%3329) ;
                                                                                                                                           mul_add[0][88]<=((mult_out_00[88] + mult_out_01[88] + mult_out_02[88])%3329) ;
                                                                                                                                           mul_add[0][89]<=((mult_out_00[89] + mult_out_01[89] + mult_out_02[89])%3329) ;
                                                                                                                                           mul_add[0][90]<=((mult_out_00[90] + mult_out_01[90] + mult_out_02[90])%3329) ;
                                                                                                                                           mul_add[0][91]<=((mult_out_00[91] + mult_out_01[91] + mult_out_02[91])%3329) ;
                                                                                                                                           mul_add[0][92]<=((mult_out_00[92] + mult_out_01[92] + mult_out_02[92])%3329) ;
                                                                                                                                           mul_add[0][93]<=((mult_out_00[93] + mult_out_01[93] + mult_out_02[93])%3329) ;
                                                                                                                                           mul_add[0][94]<=((mult_out_00[94] + mult_out_01[94] + mult_out_02[94])%3329) ;
                                                                                                                                           mul_add[0][95]<=((mult_out_00[95] + mult_out_01[95] + mult_out_02[95])%3329) ;
                                                                                                                                           mul_add[0][96]<=((mult_out_00[96] + mult_out_01[96] + mult_out_02[96])%3329) ;
                                                                                                                                           mul_add[0][97]<=((mult_out_00[97] + mult_out_01[97] + mult_out_02[97])%3329) ;
                                                                                                                                           mul_add[0][98]<=((mult_out_00[98] + mult_out_01[98] + mult_out_02[98])%3329) ;
                                                                                                                                           mul_add[0][99]<=((mult_out_00[99] + mult_out_01[99] + mult_out_02[99])%3329) ;
                                                                                                                                           mul_add[0][100]<=((mult_out_00[100] + mult_out_01[100] + mult_out_02[100])%3329) ;
                                                                                                                                           mul_add[0][101]<=((mult_out_00[101] + mult_out_01[101] + mult_out_02[101])%3329) ;
                                                                                                                                           mul_add[0][102]<=((mult_out_00[102] + mult_out_01[102] + mult_out_02[102])%3329) ;
                                                                                                                                           mul_add[0][103]<=((mult_out_00[103] + mult_out_01[103] + mult_out_02[103])%3329) ;
                                                                                                                                           mul_add[0][104]<=((mult_out_00[104] + mult_out_01[104] + mult_out_02[104])%3329) ;
                                                                                                                                           mul_add[0][105]<=((mult_out_00[105] + mult_out_01[105] + mult_out_02[105])%3329) ;
                                                                                                                                           mul_add[0][106]<=((mult_out_00[106] + mult_out_01[106] + mult_out_02[106])%3329) ;
                                                                                                                                           mul_add[0][107]<=((mult_out_00[107] + mult_out_01[107] + mult_out_02[107])%3329) ;
                                                                                                                                           mul_add[0][108]<=((mult_out_00[108] + mult_out_01[108] + mult_out_02[108])%3329) ;
                                                                                                                                           mul_add[0][109]<=((mult_out_00[109] + mult_out_01[109] + mult_out_02[109])%3329) ;
                                                                                                                                           mul_add[0][110]<=((mult_out_00[110] + mult_out_01[110] + mult_out_02[110])%3329) ;
                                                                                                                                           mul_add[0][111]<=((mult_out_00[111] + mult_out_01[111] + mult_out_02[111])%3329) ;
                                                                                                                                           mul_add[0][112]<=((mult_out_00[112] + mult_out_01[112] + mult_out_02[112])%3329) ;
                                                                                                                                           mul_add[0][113]<=((mult_out_00[113] + mult_out_01[113] + mult_out_02[113])%3329) ;
                                                                                                                                           mul_add[0][114]<=((mult_out_00[114] + mult_out_01[114] + mult_out_02[114])%3329) ;
                                                                                                                                           mul_add[0][115]<=((mult_out_00[115] + mult_out_01[115] + mult_out_02[115])%3329) ;
                                                                                                                                           mul_add[0][116]<=((mult_out_00[116] + mult_out_01[116] + mult_out_02[116])%3329) ;
                                                                                                                                           mul_add[0][117]<=((mult_out_00[117] + mult_out_01[117] + mult_out_02[117])%3329) ;
                                                                                                                                           mul_add[0][118]<=((mult_out_00[118] + mult_out_01[118] + mult_out_02[118])%3329) ;
                                                                                                                                           mul_add[0][119]<=((mult_out_00[119] + mult_out_01[119] + mult_out_02[119])%3329) ;
                                                                                                                                           mul_add[0][120]<=((mult_out_00[120] + mult_out_01[120] + mult_out_02[120])%3329) ;
                                                                                                                                           mul_add[0][121]<=((mult_out_00[121] + mult_out_01[121] + mult_out_02[121])%3329) ;
                                                                                                                                           mul_add[0][122]<=((mult_out_00[122] + mult_out_01[122] + mult_out_02[122])%3329) ;
                                                                                                                                           mul_add[0][123]<=((mult_out_00[123] + mult_out_01[123] + mult_out_02[123])%3329) ;
                                                                                                                                           mul_add[0][124]<=((mult_out_00[124] + mult_out_01[124] + mult_out_02[124])%3329) ;
                                                                                                                                           mul_add[0][125]<=((mult_out_00[125] + mult_out_01[125] + mult_out_02[125])%3329) ;
                                                                                                                                           mul_add[0][126]<=((mult_out_00[126] + mult_out_01[126] + mult_out_02[126])%3329) ;
                                                                                                                                           mul_add[0][127]<=((mult_out_00[127] + mult_out_01[127] + mult_out_02[127])%3329) ;
                                                                                                                                           mul_add[0][128]<=((mult_out_00[128] + mult_out_01[128] + mult_out_02[128])%3329) ;
                                                                                                                                           mul_add[0][129]<=((mult_out_00[129] + mult_out_01[129] + mult_out_02[129])%3329) ;
                                                                                                                                           mul_add[0][130]<=((mult_out_00[130] + mult_out_01[130] + mult_out_02[130])%3329) ;
                                                                                                                                           mul_add[0][131]<=((mult_out_00[131] + mult_out_01[131] + mult_out_02[131])%3329) ;
                                                                                                                                           mul_add[0][132]<=((mult_out_00[132] + mult_out_01[132] + mult_out_02[132])%3329) ;
                                                                                                                                           mul_add[0][133]<=((mult_out_00[133] + mult_out_01[133] + mult_out_02[133])%3329) ;
                                                                                                                                           mul_add[0][134]<=((mult_out_00[134] + mult_out_01[134] + mult_out_02[134])%3329) ;
                                                                                                                                           mul_add[0][135]<=((mult_out_00[135] + mult_out_01[135] + mult_out_02[135])%3329) ;
                                                                                                                                           mul_add[0][136]<=((mult_out_00[136] + mult_out_01[136] + mult_out_02[136])%3329) ;
                                                                                                                                           mul_add[0][137]<=((mult_out_00[137] + mult_out_01[137] + mult_out_02[137])%3329) ;
                                                                                                                                           mul_add[0][138]<=((mult_out_00[138] + mult_out_01[138] + mult_out_02[138])%3329) ;
                                                                                                                                           mul_add[0][139]<=((mult_out_00[139] + mult_out_01[139] + mult_out_02[139])%3329) ;
                                                                                                                                           mul_add[0][140]<=((mult_out_00[140] + mult_out_01[140] + mult_out_02[140])%3329) ;
                                                                                                                                           mul_add[0][141]<=((mult_out_00[141] + mult_out_01[141] + mult_out_02[141])%3329) ;
                                                                                                                                           mul_add[0][142]<=((mult_out_00[142] + mult_out_01[142] + mult_out_02[142])%3329) ;
                                                                                                                                           mul_add[0][143]<=((mult_out_00[143] + mult_out_01[143] + mult_out_02[143])%3329) ;
                                                                                                                                           mul_add[0][144]<=((mult_out_00[144] + mult_out_01[144] + mult_out_02[144])%3329) ;
                                                                                                                                           mul_add[0][145]<=((mult_out_00[145] + mult_out_01[145] + mult_out_02[145])%3329) ;
                                                                                                                                           mul_add[0][146]<=((mult_out_00[146] + mult_out_01[146] + mult_out_02[146])%3329) ;
                                                                                                                                           mul_add[0][147]<=((mult_out_00[147] + mult_out_01[147] + mult_out_02[147])%3329) ;
                                                                                                                                           mul_add[0][148]<=((mult_out_00[148] + mult_out_01[148] + mult_out_02[148])%3329) ;
                                                                                                                                           mul_add[0][149]<=((mult_out_00[149] + mult_out_01[149] + mult_out_02[149])%3329) ;
                                                                                                                                           mul_add[0][150]<=((mult_out_00[150] + mult_out_01[150] + mult_out_02[150])%3329) ;
                                                                                                                                           mul_add[0][151]<=((mult_out_00[151] + mult_out_01[151] + mult_out_02[151])%3329) ;
                                                                                                                                           mul_add[0][152]<=((mult_out_00[152] + mult_out_01[152] + mult_out_02[152])%3329) ;
                                                                                                                                           mul_add[0][153]<=((mult_out_00[153] + mult_out_01[153] + mult_out_02[153])%3329) ;
                                                                                                                                           mul_add[0][154]<=((mult_out_00[154] + mult_out_01[154] + mult_out_02[154])%3329) ;
                                                                                                                                           mul_add[0][155]<=((mult_out_00[155] + mult_out_01[155] + mult_out_02[155])%3329) ;
                                                                                                                                           mul_add[0][156]<=((mult_out_00[156] + mult_out_01[156] + mult_out_02[156])%3329) ;
                                                                                                                                           mul_add[0][157]<=((mult_out_00[157] + mult_out_01[157] + mult_out_02[157])%3329) ;
                                                                                                                                           mul_add[0][158]<=((mult_out_00[158] + mult_out_01[158] + mult_out_02[158])%3329) ;
                                                                                                                                           mul_add[0][159]<=((mult_out_00[159] + mult_out_01[159] + mult_out_02[159])%3329) ;
                                                                                                                                           mul_add[0][160]<=((mult_out_00[160] + mult_out_01[160] + mult_out_02[160])%3329) ;
                                                                                                                                           mul_add[0][161]<=((mult_out_00[161] + mult_out_01[161] + mult_out_02[161])%3329) ;
                                                                                                                                           mul_add[0][162]<=((mult_out_00[162] + mult_out_01[162] + mult_out_02[162])%3329) ;
                                                                                                                                           mul_add[0][163]<=((mult_out_00[163] + mult_out_01[163] + mult_out_02[163])%3329) ;
                                                                                                                                           mul_add[0][164]<=((mult_out_00[164] + mult_out_01[164] + mult_out_02[164])%3329) ;
                                                                                                                                           mul_add[0][165]<=((mult_out_00[165] + mult_out_01[165] + mult_out_02[165])%3329) ;
                                                                                                                                           mul_add[0][166]<=((mult_out_00[166] + mult_out_01[166] + mult_out_02[166])%3329) ;
                                                                                                                                           mul_add[0][167]<=((mult_out_00[167] + mult_out_01[167] + mult_out_02[167])%3329) ;
                                                                                                                                           mul_add[0][168]<=((mult_out_00[168] + mult_out_01[168] + mult_out_02[168])%3329) ;
                                                                                                                                           mul_add[0][169]<=((mult_out_00[169] + mult_out_01[169] + mult_out_02[169])%3329) ;
                                                                                                                                           mul_add[0][170]<=((mult_out_00[170] + mult_out_01[170] + mult_out_02[170])%3329) ;
                                                                                                                                           mul_add[0][171]<=((mult_out_00[171] + mult_out_01[171] + mult_out_02[171])%3329) ;
                                                                                                                                           mul_add[0][172]<=((mult_out_00[172] + mult_out_01[172] + mult_out_02[172])%3329) ;
                                                                                                                                           mul_add[0][173]<=((mult_out_00[173] + mult_out_01[173] + mult_out_02[173])%3329) ;
                                                                                                                                           mul_add[0][174]<=((mult_out_00[174] + mult_out_01[174] + mult_out_02[174])%3329) ;
                                                                                                                                           mul_add[0][175]<=((mult_out_00[175] + mult_out_01[175] + mult_out_02[175])%3329) ;
                                                                                                                                           mul_add[0][176]<=((mult_out_00[176] + mult_out_01[176] + mult_out_02[176])%3329) ;
                                                                                                                                           mul_add[0][177]<=((mult_out_00[177] + mult_out_01[177] + mult_out_02[177])%3329) ;
                                                                                                                                           mul_add[0][178]<=((mult_out_00[178] + mult_out_01[178] + mult_out_02[178])%3329) ;
                                                                                                                                           mul_add[0][179]<=((mult_out_00[179] + mult_out_01[179] + mult_out_02[179])%3329) ;
                                                                                                                                           mul_add[0][180]<=((mult_out_00[180] + mult_out_01[180] + mult_out_02[180])%3329) ;
                                                                                                                                           mul_add[0][181]<=((mult_out_00[181] + mult_out_01[181] + mult_out_02[181])%3329) ;
                                                                                                                                           mul_add[0][182]<=((mult_out_00[182] + mult_out_01[182] + mult_out_02[182])%3329) ;
                                                                                                                                           mul_add[0][183]<=((mult_out_00[183] + mult_out_01[183] + mult_out_02[183])%3329) ;
                                                                                                                                           mul_add[0][184]<=((mult_out_00[184] + mult_out_01[184] + mult_out_02[184])%3329) ;
                                                                                                                                           mul_add[0][185]<=((mult_out_00[185] + mult_out_01[185] + mult_out_02[185])%3329) ;
                                                                                                                                           mul_add[0][186]<=((mult_out_00[186] + mult_out_01[186] + mult_out_02[186])%3329) ;
                                                                                                                                           mul_add[0][187]<=((mult_out_00[187] + mult_out_01[187] + mult_out_02[187])%3329) ;
                                                                                                                                           mul_add[0][188]<=((mult_out_00[188] + mult_out_01[188] + mult_out_02[188])%3329) ;
                                                                                                                                           mul_add[0][189]<=((mult_out_00[189] + mult_out_01[189] + mult_out_02[189])%3329) ;
                                                                                                                                           mul_add[0][190]<=((mult_out_00[190] + mult_out_01[190] + mult_out_02[190])%3329) ;
                                                                                                                                           mul_add[0][191]<=((mult_out_00[191] + mult_out_01[191] + mult_out_02[191])%3329) ;
                                                                                                                                           mul_add[0][192]<=((mult_out_00[192] + mult_out_01[192] + mult_out_02[192])%3329) ;
                                                                                                                                           mul_add[0][193]<=((mult_out_00[193] + mult_out_01[193] + mult_out_02[193])%3329) ;
                                                                                                                                           mul_add[0][194]<=((mult_out_00[194] + mult_out_01[194] + mult_out_02[194])%3329) ;
                                                                                                                                           mul_add[0][195]<=((mult_out_00[195] + mult_out_01[195] + mult_out_02[195])%3329) ;
                                                                                                                                           mul_add[0][196]<=((mult_out_00[196] + mult_out_01[196] + mult_out_02[196])%3329) ;
                                                                                                                                           mul_add[0][197]<=((mult_out_00[197] + mult_out_01[197] + mult_out_02[197])%3329) ;
                                                                                                                                           mul_add[0][198]<=((mult_out_00[198] + mult_out_01[198] + mult_out_02[198])%3329) ;
                                                                                                                                           mul_add[0][199]<=((mult_out_00[199] + mult_out_01[199] + mult_out_02[199])%3329) ;
                                                                                                                                           mul_add[0][200]<=((mult_out_00[200] + mult_out_01[200] + mult_out_02[200])%3329) ;
                                                                                                                                           mul_add[0][201]<=((mult_out_00[201] + mult_out_01[201] + mult_out_02[201])%3329) ;
                                                                                                                                           mul_add[0][202]<=((mult_out_00[202] + mult_out_01[202] + mult_out_02[202])%3329) ;
                                                                                                                                           mul_add[0][203]<=((mult_out_00[203] + mult_out_01[203] + mult_out_02[203])%3329) ;
                                                                                                                                           mul_add[0][204]<=((mult_out_00[204] + mult_out_01[204] + mult_out_02[204])%3329) ;
                                                                                                                                           mul_add[0][205]<=((mult_out_00[205] + mult_out_01[205] + mult_out_02[205])%3329) ;
                                                                                                                                           mul_add[0][206]<=((mult_out_00[206] + mult_out_01[206] + mult_out_02[206])%3329) ;
                                                                                                                                           mul_add[0][207]<=((mult_out_00[207] + mult_out_01[207] + mult_out_02[207])%3329) ;
                                                                                                                                           mul_add[0][208]<=((mult_out_00[208] + mult_out_01[208] + mult_out_02[208])%3329) ;
                                                                                                                                           mul_add[0][209]<=((mult_out_00[209] + mult_out_01[209] + mult_out_02[209])%3329) ;
                                                                                                                                           mul_add[0][210]<=((mult_out_00[210] + mult_out_01[210] + mult_out_02[210])%3329) ;
                                                                                                                                           mul_add[0][211]<=((mult_out_00[211] + mult_out_01[211] + mult_out_02[211])%3329) ;
                                                                                                                                           mul_add[0][212]<=((mult_out_00[212] + mult_out_01[212] + mult_out_02[212])%3329) ;
                                                                                                                                           mul_add[0][213]<=((mult_out_00[213] + mult_out_01[213] + mult_out_02[213])%3329) ;
                                                                                                                                           mul_add[0][214]<=((mult_out_00[214] + mult_out_01[214] + mult_out_02[214])%3329) ;
                                                                                                                                           mul_add[0][215]<=((mult_out_00[215] + mult_out_01[215] + mult_out_02[215])%3329) ;
                                                                                                                                           mul_add[0][216]<=((mult_out_00[216] + mult_out_01[216] + mult_out_02[216])%3329) ;
                                                                                                                                           mul_add[0][217]<=((mult_out_00[217] + mult_out_01[217] + mult_out_02[217])%3329) ;
                                                                                                                                           mul_add[0][218]<=((mult_out_00[218] + mult_out_01[218] + mult_out_02[218])%3329) ;
                                                                                                                                           mul_add[0][219]<=((mult_out_00[219] + mult_out_01[219] + mult_out_02[219])%3329) ;
                                                                                                                                           mul_add[0][220]<=((mult_out_00[220] + mult_out_01[220] + mult_out_02[220])%3329) ;
                                                                                                                                           mul_add[0][221]<=((mult_out_00[221] + mult_out_01[221] + mult_out_02[221])%3329) ;
                                                                                                                                           mul_add[0][222]<=((mult_out_00[222] + mult_out_01[222] + mult_out_02[222])%3329) ;
                                                                                                                                           mul_add[0][223]<=((mult_out_00[223] + mult_out_01[223] + mult_out_02[223])%3329) ;
                                                                                                                                           mul_add[0][224]<=((mult_out_00[224] + mult_out_01[224] + mult_out_02[224])%3329) ;
                                                                                                                                           mul_add[0][225]<=((mult_out_00[225] + mult_out_01[225] + mult_out_02[225])%3329) ;
                                                                                                                                           mul_add[0][226]<=((mult_out_00[226] + mult_out_01[226] + mult_out_02[226])%3329) ;
                                                                                                                                           mul_add[0][227]<=((mult_out_00[227] + mult_out_01[227] + mult_out_02[227])%3329) ;
                                                                                                                                           mul_add[0][228]<=((mult_out_00[228] + mult_out_01[228] + mult_out_02[228])%3329) ;
                                                                                                                                           mul_add[0][229]<=((mult_out_00[229] + mult_out_01[229] + mult_out_02[229])%3329) ;
                                                                                                                                           mul_add[0][230]<=((mult_out_00[230] + mult_out_01[230] + mult_out_02[230])%3329) ;
                                                                                                                                           mul_add[0][231]<=((mult_out_00[231] + mult_out_01[231] + mult_out_02[231])%3329) ;
                                                                                                                                           mul_add[0][232]<=((mult_out_00[232] + mult_out_01[232] + mult_out_02[232])%3329) ;
                                                                                                                                           mul_add[0][233]<=((mult_out_00[233] + mult_out_01[233] + mult_out_02[233])%3329) ;
                                                                                                                                           mul_add[0][234]<=((mult_out_00[234] + mult_out_01[234] + mult_out_02[234])%3329) ;
                                                                                                                                           mul_add[0][235]<=((mult_out_00[235] + mult_out_01[235] + mult_out_02[235])%3329) ;
                                                                                                                                           mul_add[0][236]<=((mult_out_00[236] + mult_out_01[236] + mult_out_02[236])%3329) ;
                                                                                                                                           mul_add[0][237]<=((mult_out_00[237] + mult_out_01[237] + mult_out_02[237])%3329) ;
                                                                                                                                           mul_add[0][238]<=((mult_out_00[238] + mult_out_01[238] + mult_out_02[238])%3329) ;
                                                                                                                                           mul_add[0][239]<=((mult_out_00[239] + mult_out_01[239] + mult_out_02[239])%3329) ;
                                                                                                                                           mul_add[0][240]<=((mult_out_00[240] + mult_out_01[240] + mult_out_02[240])%3329) ;
                                                                                                                                           mul_add[0][241]<=((mult_out_00[241] + mult_out_01[241] + mult_out_02[241])%3329) ;
                                                                                                                                           mul_add[0][242]<=((mult_out_00[242] + mult_out_01[242] + mult_out_02[242])%3329) ;
                                                                                                                                           mul_add[0][243]<=((mult_out_00[243] + mult_out_01[243] + mult_out_02[243])%3329) ;
                                                                                                                                           mul_add[0][244]<=((mult_out_00[244] + mult_out_01[244] + mult_out_02[244])%3329) ;
                                                                                                                                           mul_add[0][245]<=((mult_out_00[245] + mult_out_01[245] + mult_out_02[245])%3329) ;
                                                                                                                                           mul_add[0][246]<=((mult_out_00[246] + mult_out_01[246] + mult_out_02[246])%3329) ;
                                                                                                                                           mul_add[0][247]<=((mult_out_00[247] + mult_out_01[247] + mult_out_02[247])%3329) ;
                                                                                                                                           mul_add[0][248]<=((mult_out_00[248] + mult_out_01[248] + mult_out_02[248])%3329) ;
                                                                                                                                           mul_add[0][249]<=((mult_out_00[249] + mult_out_01[249] + mult_out_02[249])%3329) ;
                                                                                                                                           mul_add[0][250]<=((mult_out_00[250] + mult_out_01[250] + mult_out_02[250])%3329) ;
                                                                                                                                           mul_add[0][251]<=((mult_out_00[251] + mult_out_01[251] + mult_out_02[251])%3329) ;
                                                                                                                                           mul_add[0][252]<=((mult_out_00[252] + mult_out_01[252] + mult_out_02[252])%3329) ;
                                                                                                                                           mul_add[0][253]<=((mult_out_00[253] + mult_out_01[253] + mult_out_02[253])%3329) ;
                                                                                                                                           mul_add[0][254]<=((mult_out_00[254] + mult_out_01[254] + mult_out_02[254])%3329) ;
                                                                                                                                           mul_add[0][255]<=((mult_out_00[255] + mult_out_01[255] + mult_out_02[255])%3329) ;
                                                                                                                                          
                                                                                                                                           mul_add[1][0]<=((mult_out_10[0] + mult_out_11[0] + mult_out_12[0])%3329) ;
                                                                                                                                           mul_add[1][1]<=((mult_out_10[1] + mult_out_11[1] + mult_out_12[1])%3329) ;
                                                                                                                                           mul_add[1][2]<=((mult_out_10[2] + mult_out_11[2] + mult_out_12[2])%3329) ;
                                                                                                                                           mul_add[1][3]<=((mult_out_10[3] + mult_out_11[3] + mult_out_12[3])%3329) ;
                                                                                                                                           mul_add[1][4]<=((mult_out_10[4] + mult_out_11[4] + mult_out_12[4])%3329) ;
                                                                                                                                           mul_add[1][5]<=((mult_out_10[5] + mult_out_11[5] + mult_out_12[5])%3329) ;
                                                                                                                                           mul_add[1][6]<=((mult_out_10[6] + mult_out_11[6] + mult_out_12[6])%3329) ;
                                                                                                                                           mul_add[1][7]<=((mult_out_10[7] + mult_out_11[7] + mult_out_12[7])%3329) ;
                                                                                                                                           mul_add[1][8]<=((mult_out_10[8] + mult_out_11[8] + mult_out_12[8])%3329) ;
                                                                                                                                           mul_add[1][9]<=((mult_out_10[9] + mult_out_11[9] + mult_out_12[9])%3329) ;
                                                                                                                                           mul_add[1][10]<=((mult_out_10[10] + mult_out_11[10] + mult_out_12[10])%3329) ;
                                                                                                                                           mul_add[1][11]<=((mult_out_10[11] + mult_out_11[11] + mult_out_12[11])%3329) ;
                                                                                                                                           mul_add[1][12]<=((mult_out_10[12] + mult_out_11[12] + mult_out_12[12])%3329) ;
                                                                                                                                           mul_add[1][13]<=((mult_out_10[13] + mult_out_11[13] + mult_out_12[13])%3329) ;
                                                                                                                                           mul_add[1][14]<=((mult_out_10[14] + mult_out_11[14] + mult_out_12[14])%3329) ;
                                                                                                                                           mul_add[1][15]<=((mult_out_10[15] + mult_out_11[15] + mult_out_12[15])%3329) ;
                                                                                                                                           mul_add[1][16]<=((mult_out_10[16] + mult_out_11[16] + mult_out_12[16])%3329) ;
                                                                                                                                           mul_add[1][17]<=((mult_out_10[17] + mult_out_11[17] + mult_out_12[17])%3329) ;
                                                                                                                                           mul_add[1][18]<=((mult_out_10[18] + mult_out_11[18] + mult_out_12[18])%3329) ;
                                                                                                                                           mul_add[1][19]<=((mult_out_10[19] + mult_out_11[19] + mult_out_12[19])%3329) ;
                                                                                                                                           mul_add[1][20]<=((mult_out_10[20] + mult_out_11[20] + mult_out_12[20])%3329) ;
                                                                                                                                           mul_add[1][21]<=((mult_out_10[21] + mult_out_11[21] + mult_out_12[21])%3329) ;
                                                                                                                                           mul_add[1][22]<=((mult_out_10[22] + mult_out_11[22] + mult_out_12[22])%3329) ;
                                                                                                                                           mul_add[1][23]<=((mult_out_10[23] + mult_out_11[23] + mult_out_12[23])%3329) ;
                                                                                                                                           mul_add[1][24]<=((mult_out_10[24] + mult_out_11[24] + mult_out_12[24])%3329) ;
                                                                                                                                           mul_add[1][25]<=((mult_out_10[25] + mult_out_11[25] + mult_out_12[25])%3329) ;
                                                                                                                                           mul_add[1][26]<=((mult_out_10[26] + mult_out_11[26] + mult_out_12[26])%3329) ;
                                                                                                                                           mul_add[1][27]<=((mult_out_10[27] + mult_out_11[27] + mult_out_12[27])%3329) ;
                                                                                                                                           mul_add[1][28]<=((mult_out_10[28] + mult_out_11[28] + mult_out_12[28])%3329) ;
                                                                                                                                           mul_add[1][29]<=((mult_out_10[29] + mult_out_11[29] + mult_out_12[29])%3329) ;
                                                                                                                                           mul_add[1][30]<=((mult_out_10[30] + mult_out_11[30] + mult_out_12[30])%3329) ;
                                                                                                                                           mul_add[1][31]<=((mult_out_10[31] + mult_out_11[31] + mult_out_12[31])%3329) ;
                                                                                                                                           mul_add[1][32]<=((mult_out_10[32] + mult_out_11[32] + mult_out_12[32])%3329) ;
                                                                                                                                           mul_add[1][33]<=((mult_out_10[33] + mult_out_11[33] + mult_out_12[33])%3329) ;
                                                                                                                                           mul_add[1][34]<=((mult_out_10[34] + mult_out_11[34] + mult_out_12[34])%3329) ;
                                                                                                                                           mul_add[1][35]<=((mult_out_10[35] + mult_out_11[35] + mult_out_12[35])%3329) ;
                                                                                                                                           mul_add[1][36]<=((mult_out_10[36] + mult_out_11[36] + mult_out_12[36])%3329) ;
                                                                                                                                           mul_add[1][37]<=((mult_out_10[37] + mult_out_11[37] + mult_out_12[37])%3329) ;
                                                                                                                                           mul_add[1][38]<=((mult_out_10[38] + mult_out_11[38] + mult_out_12[38])%3329) ;
                                                                                                                                           mul_add[1][39]<=((mult_out_10[39] + mult_out_11[39] + mult_out_12[39])%3329) ;
                                                                                                                                           mul_add[1][40]<=((mult_out_10[40] + mult_out_11[40] + mult_out_12[40])%3329) ;
                                                                                                                                           mul_add[1][41]<=((mult_out_10[41] + mult_out_11[41] + mult_out_12[41])%3329) ;
                                                                                                                                           mul_add[1][42]<=((mult_out_10[42] + mult_out_11[42] + mult_out_12[42])%3329) ;
                                                                                                                                           mul_add[1][43]<=((mult_out_10[43] + mult_out_11[43] + mult_out_12[43])%3329) ;
                                                                                                                                           mul_add[1][44]<=((mult_out_10[44] + mult_out_11[44] + mult_out_12[44])%3329) ;
                                                                                                                                           mul_add[1][45]<=((mult_out_10[45] + mult_out_11[45] + mult_out_12[45])%3329) ;
                                                                                                                                           mul_add[1][46]<=((mult_out_10[46] + mult_out_11[46] + mult_out_12[46])%3329) ;
                                                                                                                                           mul_add[1][47]<=((mult_out_10[47] + mult_out_11[47] + mult_out_12[47])%3329) ;
                                                                                                                                           mul_add[1][48]<=((mult_out_10[48] + mult_out_11[48] + mult_out_12[48])%3329) ;
                                                                                                                                           mul_add[1][49]<=((mult_out_10[49] + mult_out_11[49] + mult_out_12[49])%3329) ;
                                                                                                                                           mul_add[1][50]<=((mult_out_10[50] + mult_out_11[50] + mult_out_12[50])%3329) ;
                                                                                                                                           mul_add[1][51]<=((mult_out_10[51] + mult_out_11[51] + mult_out_12[51])%3329) ;
                                                                                                                                           mul_add[1][52]<=((mult_out_10[52] + mult_out_11[52] + mult_out_12[52])%3329) ;
                                                                                                                                           mul_add[1][53]<=((mult_out_10[53] + mult_out_11[53] + mult_out_12[53])%3329) ;
                                                                                                                                           mul_add[1][54]<=((mult_out_10[54] + mult_out_11[54] + mult_out_12[54])%3329) ;
                                                                                                                                           mul_add[1][55]<=((mult_out_10[55] + mult_out_11[55] + mult_out_12[55])%3329) ;
                                                                                                                                           mul_add[1][56]<=((mult_out_10[56] + mult_out_11[56] + mult_out_12[56])%3329) ;
                                                                                                                                           mul_add[1][57]<=((mult_out_10[57] + mult_out_11[57] + mult_out_12[57])%3329) ;
                                                                                                                                           mul_add[1][58]<=((mult_out_10[58] + mult_out_11[58] + mult_out_12[58])%3329) ;
                                                                                                                                           mul_add[1][59]<=((mult_out_10[59] + mult_out_11[59] + mult_out_12[59])%3329) ;
                                                                                                                                           mul_add[1][60]<=((mult_out_10[60] + mult_out_11[60] + mult_out_12[60])%3329) ;
                                                                                                                                           mul_add[1][61]<=((mult_out_10[61] + mult_out_11[61] + mult_out_12[61])%3329) ;
                                                                                                                                           mul_add[1][62]<=((mult_out_10[62] + mult_out_11[62] + mult_out_12[62])%3329) ;
                                                                                                                                           mul_add[1][63]<=((mult_out_10[63] + mult_out_11[63] + mult_out_12[63])%3329) ;
                                                                                                                                           mul_add[1][64]<=((mult_out_10[64] + mult_out_11[64] + mult_out_12[64])%3329) ;
                                                                                                                                           mul_add[1][65]<=((mult_out_10[65] + mult_out_11[65] + mult_out_12[65])%3329) ;
                                                                                                                                           mul_add[1][66]<=((mult_out_10[66] + mult_out_11[66] + mult_out_12[66])%3329) ;
                                                                                                                                           mul_add[1][67]<=((mult_out_10[67] + mult_out_11[67] + mult_out_12[67])%3329) ;
                                                                                                                                           mul_add[1][68]<=((mult_out_10[68] + mult_out_11[68] + mult_out_12[68])%3329) ;
                                                                                                                                           mul_add[1][69]<=((mult_out_10[69] + mult_out_11[69] + mult_out_12[69])%3329) ;
                                                                                                                                           mul_add[1][70]<=((mult_out_10[70] + mult_out_11[70] + mult_out_12[70])%3329) ;
                                                                                                                                           mul_add[1][71]<=((mult_out_10[71] + mult_out_11[71] + mult_out_12[71])%3329) ;
                                                                                                                                           mul_add[1][72]<=((mult_out_10[72] + mult_out_11[72] + mult_out_12[72])%3329) ;
                                                                                                                                           mul_add[1][73]<=((mult_out_10[73] + mult_out_11[73] + mult_out_12[73])%3329) ;
                                                                                                                                           mul_add[1][74]<=((mult_out_10[74] + mult_out_11[74] + mult_out_12[74])%3329) ;
                                                                                                                                           mul_add[1][75]<=((mult_out_10[75] + mult_out_11[75] + mult_out_12[75])%3329) ;
                                                                                                                                           mul_add[1][76]<=((mult_out_10[76] + mult_out_11[76] + mult_out_12[76])%3329) ;
                                                                                                                                           mul_add[1][77]<=((mult_out_10[77] + mult_out_11[77] + mult_out_12[77])%3329) ;
                                                                                                                                           mul_add[1][78]<=((mult_out_10[78] + mult_out_11[78] + mult_out_12[78])%3329) ;
                                                                                                                                           mul_add[1][79]<=((mult_out_10[79] + mult_out_11[79] + mult_out_12[79])%3329) ;
                                                                                                                                           mul_add[1][80]<=((mult_out_10[80] + mult_out_11[80] + mult_out_12[80])%3329) ;
                                                                                                                                           mul_add[1][81]<=((mult_out_10[81] + mult_out_11[81] + mult_out_12[81])%3329) ;
                                                                                                                                           mul_add[1][82]<=((mult_out_10[82] + mult_out_11[82] + mult_out_12[82])%3329) ;
                                                                                                                                           mul_add[1][83]<=((mult_out_10[83] + mult_out_11[83] + mult_out_12[83])%3329) ;
                                                                                                                                           mul_add[1][84]<=((mult_out_10[84] + mult_out_11[84] + mult_out_12[84])%3329) ;
                                                                                                                                           mul_add[1][85]<=((mult_out_10[85] + mult_out_11[85] + mult_out_12[85])%3329) ;
                                                                                                                                           mul_add[1][86]<=((mult_out_10[86] + mult_out_11[86] + mult_out_12[86])%3329) ;
                                                                                                                                           mul_add[1][87]<=((mult_out_10[87] + mult_out_11[87] + mult_out_12[87])%3329) ;
                                                                                                                                           mul_add[1][88]<=((mult_out_10[88] + mult_out_11[88] + mult_out_12[88])%3329) ;
                                                                                                                                           mul_add[1][89]<=((mult_out_10[89] + mult_out_11[89] + mult_out_12[89])%3329) ;
                                                                                                                                           mul_add[1][90]<=((mult_out_10[90] + mult_out_11[90] + mult_out_12[90])%3329) ;
                                                                                                                                           mul_add[1][91]<=((mult_out_10[91] + mult_out_11[91] + mult_out_12[91])%3329) ;
                                                                                                                                           mul_add[1][92]<=((mult_out_10[92] + mult_out_11[92] + mult_out_12[92])%3329) ;
                                                                                                                                           mul_add[1][93]<=((mult_out_10[93] + mult_out_11[93] + mult_out_12[93])%3329) ;
                                                                                                                                           mul_add[1][94]<=((mult_out_10[94] + mult_out_11[94] + mult_out_12[94])%3329) ;
                                                                                                                                           mul_add[1][95]<=((mult_out_10[95] + mult_out_11[95] + mult_out_12[95])%3329) ;
                                                                                                                                           mul_add[1][96]<=((mult_out_10[96] + mult_out_11[96] + mult_out_12[96])%3329) ;
                                                                                                                                           mul_add[1][97]<=((mult_out_10[97] + mult_out_11[97] + mult_out_12[97])%3329) ;
                                                                                                                                           mul_add[1][98]<=((mult_out_10[98] + mult_out_11[98] + mult_out_12[98])%3329) ;
                                                                                                                                           mul_add[1][99]<=((mult_out_10[99] + mult_out_11[99] + mult_out_12[99])%3329) ;
                                                                                                                                           mul_add[1][100]<=((mult_out_10[100] + mult_out_11[100] + mult_out_12[100])%3329);
                                                                                                                                           mul_add[1][101]<=((mult_out_10[101] + mult_out_11[101] + mult_out_12[101])%3329) ;
                                                                                                                                           mul_add[1][102]<=((mult_out_10[102] + mult_out_11[102] + mult_out_12[102])%3329) ;
                                                                                                                                           mul_add[1][103]<=((mult_out_10[103] + mult_out_11[103] + mult_out_12[103])%3329) ;
                                                                                                                                           mul_add[1][104]<=((mult_out_10[104] + mult_out_11[104] + mult_out_12[104])%3329) ;
                                                                                                                                           mul_add[1][105]<=((mult_out_10[105] + mult_out_11[105] + mult_out_12[105])%3329) ;
                                                                                                                                           mul_add[1][106]<=((mult_out_10[106] + mult_out_11[106] + mult_out_12[106])%3329) ;
                                                                                                                                           mul_add[1][107]<=((mult_out_10[107] + mult_out_11[107] + mult_out_12[107])%3329) ;
                                                                                                                                           mul_add[1][108]<=((mult_out_10[108] + mult_out_11[108] + mult_out_12[108])%3329) ;
                                                                                                                                           mul_add[1][109]<=((mult_out_10[109] + mult_out_11[109] + mult_out_12[109])%3329) ;
                                                                                                                                           mul_add[1][110]<=((mult_out_10[110] + mult_out_11[110] + mult_out_12[110])%3329) ;
                                                                                                                                           mul_add[1][111]<=((mult_out_10[111] + mult_out_11[111] + mult_out_12[111])%3329) ;
                                                                                                                                           mul_add[1][112]<=((mult_out_10[112] + mult_out_11[112] + mult_out_12[112])%3329) ;
                                                                                                                                           mul_add[1][113]<=((mult_out_10[113] + mult_out_11[113] + mult_out_12[113])%3329) ;
                                                                                                                                           mul_add[1][114]<=((mult_out_10[114] + mult_out_11[114] + mult_out_12[114])%3329) ;
                                                                                                                                           mul_add[1][115]<=((mult_out_10[115] + mult_out_11[115] + mult_out_12[115])%3329) ;
                                                                                                                                           mul_add[1][116]<=((mult_out_10[116] + mult_out_11[116] + mult_out_12[116])%3329) ;
                                                                                                                                           mul_add[1][117]<=((mult_out_10[117] + mult_out_11[117] + mult_out_12[117])%3329) ;
                                                                                                                                           mul_add[1][118]<=((mult_out_10[118] + mult_out_11[118] + mult_out_12[118])%3329) ;
                                                                                                                                           mul_add[1][119]<=((mult_out_10[119] + mult_out_11[119] + mult_out_12[119])%3329) ;
                                                                                                                                           mul_add[1][120]<=((mult_out_10[120] + mult_out_11[120] + mult_out_12[120])%3329) ;
                                                                                                                                           mul_add[1][121]<=((mult_out_10[121] + mult_out_11[121] + mult_out_12[121])%3329) ;
                                                                                                                                           mul_add[1][122]<=((mult_out_10[122] + mult_out_11[122] + mult_out_12[122])%3329) ;
                                                                                                                                           mul_add[1][123]<=((mult_out_10[123] + mult_out_11[123] + mult_out_12[123])%3329);
                                                                                                                                           mul_add[1][124]<=((mult_out_10[124] + mult_out_11[124] + mult_out_12[124])%3329);
                                                                                                                                           mul_add[1][125]<=((mult_out_10[125] + mult_out_11[125] + mult_out_12[125])%3329);
                                                                                                                                           mul_add[1][126]<=((mult_out_10[126] + mult_out_11[126] + mult_out_12[126])%3329);
                                                                                                                                           mul_add[1][127]<=((mult_out_10[127] + mult_out_11[127] + mult_out_12[127])%3329);
                                                                                                                                           mul_add[1][128]<=((mult_out_10[128] + mult_out_11[128] + mult_out_12[128])%3329);
                                                                                                                                           mul_add[1][129]<=((mult_out_10[129] + mult_out_11[129] + mult_out_12[129])%3329);
                                                                                                                                           mul_add[1][130]<=((mult_out_10[130] + mult_out_11[130] + mult_out_12[130])%3329);
                                                                                                                                           mul_add[1][131]<=((mult_out_10[131] + mult_out_11[131] + mult_out_12[131])%3329);
                                                                                                                                           mul_add[1][132]<=((mult_out_10[132] + mult_out_11[132] + mult_out_12[132])%3329);
                                                                                                                                           mul_add[1][133]<=((mult_out_10[133] + mult_out_11[133] + mult_out_12[133])%3329);
                                                                                                                                           mul_add[1][134]<=((mult_out_10[134] + mult_out_11[134] + mult_out_12[134])%3329);
                                                                                                                                           mul_add[1][135]<=((mult_out_10[135] + mult_out_11[135] + mult_out_12[135])%3329);
                                                                                                                                           mul_add[1][136]<=((mult_out_10[136] + mult_out_11[136] + mult_out_12[136])%3329);
                                                                                                                                           mul_add[1][137]<=((mult_out_10[137] + mult_out_11[137] + mult_out_12[137])%3329);
                                                                                                                                           mul_add[1][138]<=((mult_out_10[138] + mult_out_11[138] + mult_out_12[138])%3329);
                                                                                                                                           mul_add[1][139]<=((mult_out_10[139] + mult_out_11[139] + mult_out_12[139])%3329);
                                                                                                                                           mul_add[1][140]<=((mult_out_10[140] + mult_out_11[140] + mult_out_12[140])%3329);
                                                                                                                                           mul_add[1][141]<=((mult_out_10[141] + mult_out_11[141] + mult_out_12[141])%3329);
                                                                                                                                           mul_add[1][142]<=((mult_out_10[142] + mult_out_11[142] + mult_out_12[142])%3329);
                                                                                                                                           mul_add[1][143]<=((mult_out_10[143] + mult_out_11[143] + mult_out_12[143])%3329);
                                                                                                                                           mul_add[1][144]<=((mult_out_10[144] + mult_out_11[144] + mult_out_12[144])%3329);
                                                                                                                                           mul_add[1][145]<=((mult_out_10[145] + mult_out_11[145] + mult_out_12[145])%3329);
                                                                                                                                           mul_add[1][146]<=((mult_out_10[146] + mult_out_11[146] + mult_out_12[146])%3329);
                                                                                                                                           mul_add[1][147]<=((mult_out_10[147] + mult_out_11[147] + mult_out_12[147])%3329);
                                                                                                                                           mul_add[1][148]<=((mult_out_10[148] + mult_out_11[148] + mult_out_12[148])%3329);
                                                                                                                                           mul_add[1][149]<=((mult_out_10[149] + mult_out_11[149] + mult_out_12[149])%3329);
                                                                                                                                           mul_add[1][150]<=((mult_out_10[150] + mult_out_11[150] + mult_out_12[150])%3329);
                                                                                                                                           mul_add[1][151]<=((mult_out_10[151] + mult_out_11[151] + mult_out_12[151])%3329);
                                                                                                                                           mul_add[1][152]<=((mult_out_10[152] + mult_out_11[152] + mult_out_12[152])%3329);
                                                                                                                                           mul_add[1][153]<=((mult_out_10[153] + mult_out_11[153] + mult_out_12[153])%3329);
                                                                                                                                           mul_add[1][154]<=((mult_out_10[154] + mult_out_11[154] + mult_out_12[154])%3329);
                                                                                                                                           mul_add[1][155]<=((mult_out_10[155] + mult_out_11[155] + mult_out_12[155])%3329);
                                                                                                                                           mul_add[1][156]<=((mult_out_10[156] + mult_out_11[156] + mult_out_12[156])%3329);
                                                                                                                                           mul_add[1][157]<=((mult_out_10[157] + mult_out_11[157] + mult_out_12[157])%3329) ;
                                                                                                                                           mul_add[1][158]<=((mult_out_10[158] + mult_out_11[158] + mult_out_12[158])%3329) ;
                                                                                                                                           mul_add[1][159]<=((mult_out_10[159] + mult_out_11[159] + mult_out_12[159])%3329);
                                                                                                                                           mul_add[1][160]<=((mult_out_10[160] + mult_out_11[160] + mult_out_12[160])%3329) ;
                                                                                                                                           mul_add[1][161]<=((mult_out_10[161] + mult_out_11[161] + mult_out_12[161])%3329) ;
                                                                                                                                           mul_add[1][162]<=((mult_out_10[162] + mult_out_11[162] + mult_out_12[162])%3329) ;
                                                                                                                                           mul_add[1][163]<=((mult_out_10[163] + mult_out_11[163] + mult_out_12[163])%3329);
                                                                                                                                           mul_add[1][164]<=((mult_out_10[164] + mult_out_11[164] + mult_out_12[164])%3329);
                                                                                                                                           mul_add[1][165]<=((mult_out_10[165] + mult_out_11[165] + mult_out_12[165])%3329) ;
                                                                                                                                           mul_add[1][166]<=((mult_out_10[166] + mult_out_11[166] + mult_out_12[166])%3329) ;
                                                                                                                                           mul_add[1][167]<=((mult_out_10[167] + mult_out_11[167] + mult_out_12[167])%3329) ;
                                                                                                                                           mul_add[1][168]<=((mult_out_10[168] + mult_out_11[168] + mult_out_12[168])%3329) ;
                                                                                                                                           mul_add[1][169]<=((mult_out_10[169] + mult_out_11[169] + mult_out_12[169])%3329) ;
                                                                                                                                           mul_add[1][170]<=((mult_out_10[170] + mult_out_11[170] + mult_out_12[170])%3329) ;
                                                                                                                                           mul_add[1][171]<=((mult_out_10[171] + mult_out_11[171] + mult_out_12[171])%3329) ;
                                                                                                                                           mul_add[1][172]<=((mult_out_10[172] + mult_out_11[172] + mult_out_12[172])%3329) ;
                                                                                                                                           mul_add[1][173]<=((mult_out_10[173] + mult_out_11[173] + mult_out_12[173])%3329) ;
                                                                                                                                           mul_add[1][174]<=((mult_out_10[174] + mult_out_11[174] + mult_out_12[174])%3329) ;
                                                                                                                                           mul_add[1][175]<=((mult_out_10[175] + mult_out_11[175] + mult_out_12[175])%3329) ;
                                                                                                                                           mul_add[1][176]<=((mult_out_10[176] + mult_out_11[176] + mult_out_12[176])%3329) ;
                                                                                                                                           mul_add[1][177]<=((mult_out_10[177] + mult_out_11[177] + mult_out_12[177])%3329) ;
                                                                                                                                           mul_add[1][178]<=((mult_out_10[178] + mult_out_11[178] + mult_out_12[178])%3329) ;
                                                                                                                                           mul_add[1][179]<=((mult_out_10[179] + mult_out_11[179] + mult_out_12[179])%3329) ;
                                                                                                                                           mul_add[1][180]<=((mult_out_10[180] + mult_out_11[180] + mult_out_12[180])%3329) ;
                                                                                                                                           mul_add[1][181]<=((mult_out_10[181] + mult_out_11[181] + mult_out_12[181])%3329) ;
                                                                                                                                           mul_add[1][182]<=((mult_out_10[182] + mult_out_11[182] + mult_out_12[182])%3329) ;
                                                                                                                                           mul_add[1][183]<=((mult_out_10[183] + mult_out_11[183] + mult_out_12[183])%3329) ;
                                                                                                                                           mul_add[1][184]<=((mult_out_10[184] + mult_out_11[184] + mult_out_12[184])%3329) ;
                                                                                                                                           mul_add[1][185]<=((mult_out_10[185] + mult_out_11[185] + mult_out_12[185])%3329) ;
                                                                                                                                           mul_add[1][186]<=((mult_out_10[186] + mult_out_11[186] + mult_out_12[186])%3329) ;
                                                                                                                                           mul_add[1][187]<=((mult_out_10[187] + mult_out_11[187] + mult_out_12[187])%3329) ;
                                                                                                                                           mul_add[1][188]<=((mult_out_10[188] + mult_out_11[188] + mult_out_12[188])%3329) ;
                                                                                                                                           mul_add[1][189]<=((mult_out_10[189] + mult_out_11[189] + mult_out_12[189])%3329) ;
                                                                                                                                           mul_add[1][190]<=((mult_out_10[190] + mult_out_11[190] + mult_out_12[190])%3329) ;
                                                                                                                                           mul_add[1][191]<=((mult_out_10[191] + mult_out_11[191] + mult_out_12[191])%3329) ;
                                                                                                                                           mul_add[1][192]<=((mult_out_10[192] + mult_out_11[192] + mult_out_12[192])%3329) ;
                                                                                                                                           mul_add[1][193]<=((mult_out_10[193] + mult_out_11[193] + mult_out_12[193])%3329) ;
                                                                                                                                           mul_add[1][194]<=((mult_out_10[194] + mult_out_11[194] + mult_out_12[194])%3329) ;
                                                                                                                                           mul_add[1][195]<=((mult_out_10[195] + mult_out_11[195] + mult_out_12[195])%3329) ;
                                                                                                                                           mul_add[1][196]<=((mult_out_10[196] + mult_out_11[196] + mult_out_12[196])%3329) ;
                                                                                                                                           mul_add[1][197]<=((mult_out_10[197] + mult_out_11[197] + mult_out_12[197])%3329) ;
                                                                                                                                           mul_add[1][198]<=((mult_out_10[198] + mult_out_11[198] + mult_out_12[198])%3329) ;
                                                                                                                                           mul_add[1][199]<=((mult_out_10[199] + mult_out_11[199] + mult_out_12[199])%3329) ;
                                                                                                                                           mul_add[1][200]<=((mult_out_10[200] + mult_out_11[200] + mult_out_12[200])%3329) ;
                                                                                                                                           mul_add[1][201]<=((mult_out_10[201] + mult_out_11[201] + mult_out_12[201])%3329) ;
                                                                                                                                           mul_add[1][202]<=((mult_out_10[202] + mult_out_11[202] + mult_out_12[202])%3329) ;
                                                                                                                                           mul_add[1][203]<=((mult_out_10[203] + mult_out_11[203] + mult_out_12[203])%3329) ;
                                                                                                                                           mul_add[1][204]<=((mult_out_10[204] + mult_out_11[204] + mult_out_12[204])%3329) ;
                                                                                                                                           mul_add[1][205]<=((mult_out_10[205] + mult_out_11[205] + mult_out_12[205])%3329) ;
                                                                                                                                           mul_add[1][206]<=((mult_out_10[206] + mult_out_11[206] + mult_out_12[206])%3329) ;
                                                                                                                                           mul_add[1][207]<=((mult_out_10[207] + mult_out_11[207] + mult_out_12[207])%3329) ;
                                                                                                                                           mul_add[1][208]<=((mult_out_10[208] + mult_out_11[208] + mult_out_12[208])%3329) ;
                                                                                                                                           mul_add[1][209]<=((mult_out_10[209] + mult_out_11[209] + mult_out_12[209])%3329) ;
                                                                                                                                           mul_add[1][210]<=((mult_out_10[210] + mult_out_11[210] + mult_out_12[210])%3329) ;
                                                                                                                                           mul_add[1][211]<=((mult_out_10[211] + mult_out_11[211] + mult_out_12[211])%3329) ;
                                                                                                                                           mul_add[1][212]<=((mult_out_10[212] + mult_out_11[212] + mult_out_12[212])%3329) ;
                                                                                                                                           mul_add[1][213]<=((mult_out_10[213] + mult_out_11[213] + mult_out_12[213])%3329) ;
                                                                                                                                           mul_add[1][214]<=((mult_out_10[214] + mult_out_11[214] + mult_out_12[214])%3329) ;
                                                                                                                                           mul_add[1][215]<=((mult_out_10[215] + mult_out_11[215] + mult_out_12[215])%3329) ;
                                                                                                                                           mul_add[1][216]<=((mult_out_10[216] + mult_out_11[216] + mult_out_12[216])%3329) ;
                                                                                                                                           mul_add[1][217]<=((mult_out_10[217] + mult_out_11[217] + mult_out_12[217])%3329) ;
                                                                                                                                           mul_add[1][218]<=((mult_out_10[218] + mult_out_11[218] + mult_out_12[218])%3329) ;
                                                                                                                                           mul_add[1][219]<=((mult_out_10[219] + mult_out_11[219] + mult_out_12[219])%3329) ;
                                                                                                                                           mul_add[1][220]<=((mult_out_10[220] + mult_out_11[220] + mult_out_12[220])%3329) ;
                                                                                                                                           mul_add[1][221]<=((mult_out_10[221] + mult_out_11[221] + mult_out_12[221])%3329) ;
                                                                                                                                           mul_add[1][222]<=((mult_out_10[222] + mult_out_11[222] + mult_out_12[222])%3329) ;
                                                                                                                                           mul_add[1][223]<=((mult_out_10[223] + mult_out_11[223] + mult_out_12[223])%3329) ;
                                                                                                                                           mul_add[1][224]<=((mult_out_10[224] + mult_out_11[224] + mult_out_12[224])%3329) ;
                                                                                                                                           mul_add[1][225]<=((mult_out_10[225] + mult_out_11[225] + mult_out_12[225])%3329) ;
                                                                                                                                           mul_add[1][226]<=((mult_out_10[226] + mult_out_11[226] + mult_out_12[226])%3329) ;
                                                                                                                                           mul_add[1][227]<=((mult_out_10[227] + mult_out_11[227] + mult_out_12[227])%3329) ;
                                                                                                                                           mul_add[1][228]<=((mult_out_10[228] + mult_out_11[228] + mult_out_12[228])%3329) ;
                                                                                                                                           mul_add[1][229]<=((mult_out_10[229] + mult_out_11[229] + mult_out_12[229])%3329) ;
                                                                                                                                           mul_add[1][230]<=((mult_out_10[230] + mult_out_11[230] + mult_out_12[230])%3329) ;
                                                                                                                                           mul_add[1][231]<=((mult_out_10[231] + mult_out_11[231] + mult_out_12[231])%3329) ;
                                                                                                                                           mul_add[1][232]<=((mult_out_10[232] + mult_out_11[232] + mult_out_12[232])%3329) ;
                                                                                                                                           mul_add[1][233]<=((mult_out_10[233] + mult_out_11[233] + mult_out_12[233])%3329) ;
                                                                                                                                           mul_add[1][234]<=((mult_out_10[234] + mult_out_11[234] + mult_out_12[234])%3329) ;
                                                                                                                                           mul_add[1][235]<=((mult_out_10[235] + mult_out_11[235] + mult_out_12[235])%3329) ;
                                                                                                                                           mul_add[1][236]<=((mult_out_10[236] + mult_out_11[236] + mult_out_12[236])%3329) ;
                                                                                                                                           mul_add[1][237]<=((mult_out_10[237] + mult_out_11[237] + mult_out_12[237])%3329) ;
                                                                                                                                           mul_add[1][238]<=((mult_out_10[238] + mult_out_11[238] + mult_out_12[238])%3329) ;
                                                                                                                                           mul_add[1][239]<=((mult_out_10[239] + mult_out_11[239] + mult_out_12[239])%3329) ;
                                                                                                                                           mul_add[1][240]<=((mult_out_10[240] + mult_out_11[240] + mult_out_12[240])%3329) ;
                                                                                                                                           mul_add[1][241]<=((mult_out_10[241] + mult_out_11[241] + mult_out_12[241])%3329) ;
                                                                                                                                           mul_add[1][242]<=((mult_out_10[242] + mult_out_11[242] + mult_out_12[242])%3329) ;
                                                                                                                                           mul_add[1][243]<=((mult_out_10[243] + mult_out_11[243] + mult_out_12[243])%3329) ;
                                                                                                                                           mul_add[1][244]<=((mult_out_10[244] + mult_out_11[244] + mult_out_12[244])%3329) ;
                                                                                                                                           mul_add[1][245]<=((mult_out_10[245] + mult_out_11[245] + mult_out_12[245])%3329) ;
                                                                                                                                           mul_add[1][246]<=((mult_out_10[246] + mult_out_11[246] + mult_out_12[246])%3329) ;
                                                                                                                                           mul_add[1][247]<=((mult_out_10[247] + mult_out_11[247] + mult_out_12[247])%3329);
                                                                                                                                           mul_add[1][248]<=((mult_out_10[248] + mult_out_11[248] + mult_out_12[248])%3329) ;
                                                                                                                                           mul_add[1][249]<=((mult_out_10[249] + mult_out_11[249] + mult_out_12[249])%3329) ;
                                                                                                                                           mul_add[1][250]<=((mult_out_10[250] + mult_out_11[250] + mult_out_12[250])%3329) ;
                                                                                                                                           mul_add[1][251]<=((mult_out_10[251] + mult_out_11[251] + mult_out_12[251])%3329) ;
                                                                                                                                           mul_add[1][252]<=((mult_out_10[252] + mult_out_11[252] + mult_out_12[252])%3329) ;
                                                                                                                                           mul_add[1][253]<=((mult_out_10[253] + mult_out_11[253] + mult_out_12[253])%3329) ;
                                                                                                                                           mul_add[1][254]<=((mult_out_10[254] + mult_out_11[254] + mult_out_12[254])%3329) ;
                                                                                                                                           mul_add[1][255]<=((mult_out_10[255] + mult_out_11[255] + mult_out_12[255])%3329) ;
                                                                                                                                          
                                                                                                                                      
                                                                                                                                           mul_add[2][0]<=((mult_out_20[0] + mult_out_21[0] + mult_out_22[0])%3329) ;
                                                                                                                                       mul_add[2][1]<=((mult_out_20[1] + mult_out_21[1] + mult_out_22[1])%3329) ;
                                                                                                                                       mul_add[2][2]<=((mult_out_20[2] + mult_out_21[2] + mult_out_22[2])%3329) ;
                                                                                                                                       mul_add[2][3]<=((mult_out_20[3] + mult_out_21[3] + mult_out_22[3])%3329) ;
                                                                                                                                       mul_add[2][4]<=((mult_out_20[4] + mult_out_21[4] + mult_out_22[4])%3329) ;
                                                                                                                                       mul_add[2][5]<=((mult_out_20[5] + mult_out_21[5] + mult_out_22[5])%3329) ;
                                                                                                                                       mul_add[2][6]<=((mult_out_20[6] + mult_out_21[6] + mult_out_22[6])%3329) ;
                                                                                                                                       mul_add[2][7]<=((mult_out_20[7] + mult_out_21[7] + mult_out_22[7])%3329) ;
                                                                                                                                       mul_add[2][8]<=((mult_out_20[8] + mult_out_21[8] + mult_out_22[8])%3329) ;
                                                                                                                                       mul_add[2][9]<=((mult_out_20[9] + mult_out_21[9] + mult_out_22[9])%3329) ;
                                                                                                                                       mul_add[2][10]<=((mult_out_20[10] + mult_out_21[10] + mult_out_22[10])%3329) ;
                                                                                                                                       mul_add[2][11]<=((mult_out_20[11] + mult_out_21[11] + mult_out_22[11])%3329) ;
                                                                                                                                       mul_add[2][12]<=((mult_out_20[12] + mult_out_21[12] + mult_out_22[12])%3329) ;
                                                                                                                                       mul_add[2][13]<=((mult_out_20[13] + mult_out_21[13] + mult_out_22[13])%3329) ;
                                                                                                                                       mul_add[2][14]<=((mult_out_20[14] + mult_out_21[14] + mult_out_22[14])%3329) ;
                                                                                                                                       mul_add[2][15]<=((mult_out_20[15] + mult_out_21[15] + mult_out_22[15])%3329) ;
                                                                                                                                       mul_add[2][16]<=((mult_out_20[16] + mult_out_21[16] + mult_out_22[16])%3329) ;
                                                                                                                                       mul_add[2][17]<=((mult_out_20[17] + mult_out_21[17] + mult_out_22[17])%3329) ;
                                                                                                                                       mul_add[2][18]<=((mult_out_20[18] + mult_out_21[18] + mult_out_22[18])%3329) ;
                                                                                                                                       mul_add[2][19]<=((mult_out_20[19] + mult_out_21[19] + mult_out_22[19])%3329) ;
                                                                                                                                       mul_add[2][20]<=((mult_out_20[20] + mult_out_21[20] + mult_out_22[20])%3329) ;
                                                                                                                                       mul_add[2][21]<=((mult_out_20[21] + mult_out_21[21] + mult_out_22[21])%3329) ;
                                                                                                                                       mul_add[2][22]<=((mult_out_20[22] + mult_out_21[22] + mult_out_22[22])%3329) ;
                                                                                                                                       mul_add[2][23]<=((mult_out_20[23] + mult_out_21[23] + mult_out_22[23])%3329) ;
                                                                                                                                       mul_add[2][24]<=((mult_out_20[24] + mult_out_21[24] + mult_out_22[24])%3329) ;
                                                                                                                                       mul_add[2][25]<=((mult_out_20[25] + mult_out_21[25] + mult_out_22[25])%3329) ;
                                                                                                                                       mul_add[2][26]<=((mult_out_20[26] + mult_out_21[26] + mult_out_22[26])%3329) ;
                                                                                                                                       mul_add[2][27]<=((mult_out_20[27] + mult_out_21[27] + mult_out_22[27])%3329) ;
                                                                                                                                       mul_add[2][28]<=((mult_out_20[28] + mult_out_21[28] + mult_out_22[28])%3329) ;
                                                                                                                                       mul_add[2][29]<=((mult_out_20[29] + mult_out_21[29] + mult_out_22[29])%3329) ;
                                                                                                                                       mul_add[2][30]<=((mult_out_20[30] + mult_out_21[30] + mult_out_22[30])%3329) ;
                                                                                                                                       mul_add[2][31]<=((mult_out_20[31] + mult_out_21[31] + mult_out_22[31])%3329) ;
                                                                                                                                       mul_add[2][32]<=((mult_out_20[32] + mult_out_21[32] + mult_out_22[32])%3329) ;
                                                                                                                                       mul_add[2][33]<=((mult_out_20[33] + mult_out_21[33] + mult_out_22[33])%3329) ;
                                                                                                                                       mul_add[2][34]<=((mult_out_20[34] + mult_out_21[34] + mult_out_22[34])%3329) ;
                                                                                                                                       mul_add[2][35]<=((mult_out_20[35] + mult_out_21[35] + mult_out_22[35])%3329) ;
                                                                                                                                       mul_add[2][36]<=((mult_out_20[36] + mult_out_21[36] + mult_out_22[36])%3329) ;
                                                                                                                                       mul_add[2][37]<=((mult_out_20[37] + mult_out_21[37] + mult_out_22[37])%3329) ;
                                                                                                                                       mul_add[2][38]<=((mult_out_20[38] + mult_out_21[38] + mult_out_22[38])%3329) ;
                                                                                                                                       mul_add[2][39]<=((mult_out_20[39] + mult_out_21[39] + mult_out_22[39])%3329) ;
                                                                                                                                       mul_add[2][40]<=((mult_out_20[40] + mult_out_21[40] + mult_out_22[40])%3329) ;
                                                                                                                                       mul_add[2][41]<=((mult_out_20[41] + mult_out_21[41] + mult_out_22[41])%3329) ;
                                                                                                                                       mul_add[2][42]<=((mult_out_20[42] + mult_out_21[42] + mult_out_22[42])%3329) ;
                                                                                                                                       mul_add[2][43]<=((mult_out_20[43] + mult_out_21[43] + mult_out_22[43])%3329) ;
                                                                                                                                       mul_add[2][44]<=((mult_out_20[44] + mult_out_21[44] + mult_out_22[44])%3329) ;
                                                                                                                                       mul_add[2][45]<=((mult_out_20[45] + mult_out_21[45] + mult_out_22[45])%3329) ;
                                                                                                                                       mul_add[2][46]<=((mult_out_20[46] + mult_out_21[46] + mult_out_22[46])%3329) ;
                                                                                                                                       mul_add[2][47]<=((mult_out_20[47] + mult_out_21[47] + mult_out_22[47])%3329) ;
                                                                                                                                       mul_add[2][48]<=((mult_out_20[48] + mult_out_21[48] + mult_out_22[48])%3329) ;
                                                                                                                                       mul_add[2][49]<=((mult_out_20[49] + mult_out_21[49] + mult_out_22[49])%3329) ;
                                                                                                                                       mul_add[2][50]<=((mult_out_20[50] + mult_out_21[50] + mult_out_22[50])%3329) ;
                                                                                                                                       mul_add[2][51]<=((mult_out_20[51] + mult_out_21[51] + mult_out_22[51])%3329) ;
                                                                                                                                       mul_add[2][52]<=((mult_out_20[52] + mult_out_21[52] + mult_out_22[52])%3329) ;
                                                                                                                                       mul_add[2][53]<=((mult_out_20[53] + mult_out_21[53] + mult_out_22[53])%3329) ;
                                                                                                                                       mul_add[2][54]<=((mult_out_20[54] + mult_out_21[54] + mult_out_22[54])%3329) ;
                                                                                                                                       mul_add[2][55]<=((mult_out_20[55] + mult_out_21[55] + mult_out_22[55])%3329) ;
                                                                                                                                       mul_add[2][56]<=((mult_out_20[56] + mult_out_21[56] + mult_out_22[56])%3329) ;
                                                                                                                                       mul_add[2][57]<=((mult_out_20[57] + mult_out_21[57] + mult_out_22[57])%3329) ;
                                                                                                                                       mul_add[2][58]<=((mult_out_20[58] + mult_out_21[58] + mult_out_22[58])%3329) ;
                                                                                                                                       mul_add[2][59]<=((mult_out_20[59] + mult_out_21[59] + mult_out_22[59])%3329) ;
                                                                                                                                       mul_add[2][60]<=((mult_out_20[60] + mult_out_21[60] + mult_out_22[60])%3329) ;
                                                                                                                                       mul_add[2][61]<=((mult_out_20[61] + mult_out_21[61] + mult_out_22[61])%3329) ;
                                                                                                                                       mul_add[2][62]<=((mult_out_20[62] + mult_out_21[62] + mult_out_22[62])%3329) ;
                                                                                                                                       mul_add[2][63]<=((mult_out_20[63] + mult_out_21[63] + mult_out_22[63])%3329) ;
                                                                                                                                       mul_add[2][64]<=((mult_out_20[64] + mult_out_21[64] + mult_out_22[64])%3329) ;
                                                                                                                                       mul_add[2][65]<=((mult_out_20[65] + mult_out_21[65] + mult_out_22[65])%3329) ;
                                                                                                                                       mul_add[2][66]<=((mult_out_20[66] + mult_out_21[66] + mult_out_22[66])%3329) ;
                                                                                                                                       mul_add[2][67]<=((mult_out_20[67] + mult_out_21[67] + mult_out_22[67])%3329) ;
                                                                                                                                       mul_add[2][68]<=((mult_out_20[68] + mult_out_21[68] + mult_out_22[68])%3329) ;
                                                                                                                                       mul_add[2][69]<=((mult_out_20[69] + mult_out_21[69] + mult_out_22[69])%3329) ;
                                                                                                                                       mul_add[2][70]<=((mult_out_20[70] + mult_out_21[70] + mult_out_22[70])%3329) ;
                                                                                                                                       mul_add[2][71]<=((mult_out_20[71] + mult_out_21[71] + mult_out_22[71])%3329) ;
                                                                                                                                       mul_add[2][72]<=((mult_out_20[72] + mult_out_21[72] + mult_out_22[72])%3329) ;
                                                                                                                                       mul_add[2][73]<=((mult_out_20[73] + mult_out_21[73] + mult_out_22[73])%3329) ;
                                                                                                                                       mul_add[2][74]<=((mult_out_20[74] + mult_out_21[74] + mult_out_22[74])%3329) ;
                                                                                                                                       mul_add[2][75]<=((mult_out_20[75] + mult_out_21[75] + mult_out_22[75])%3329) ;
                                                                                                                                       mul_add[2][76]<=((mult_out_20[76] + mult_out_21[76] + mult_out_22[76])%3329) ;
                                                                                                                                       mul_add[2][77]<=((mult_out_20[77] + mult_out_21[77] + mult_out_22[77])%3329) ;
                                                                                                                                       mul_add[2][78]<=((mult_out_20[78] + mult_out_21[78] + mult_out_22[78])%3329) ;
                                                                                                                                       mul_add[2][79]<=((mult_out_20[79] + mult_out_21[79] + mult_out_22[79])%3329) ;
                                                                                                                                       mul_add[2][80]<=((mult_out_20[80] + mult_out_21[80] + mult_out_22[80])%3329) ;
                                                                                                                                       mul_add[2][81]<=((mult_out_20[81] + mult_out_21[81] + mult_out_22[81])%3329) ;
                                                                                                                                       mul_add[2][82]<=((mult_out_20[82] + mult_out_21[82] + mult_out_22[82])%3329) ;
                                                                                                                                       mul_add[2][83]<=((mult_out_20[83] + mult_out_21[83] + mult_out_22[83])%3329) ;
                                                                                                                                       mul_add[2][84]<=((mult_out_20[84] + mult_out_21[84] + mult_out_22[84])%3329) ;
                                                                                                                                       mul_add[2][85]<=((mult_out_20[85] + mult_out_21[85] + mult_out_22[85])%3329) ;
                                                                                                                                       mul_add[2][86]<=((mult_out_20[86] + mult_out_21[86] + mult_out_22[86])%3329) ;
                                                                                                                                       mul_add[2][87]<=((mult_out_20[87] + mult_out_21[87] + mult_out_22[87])%3329) ;
                                                                                                                                       mul_add[2][88]<=((mult_out_20[88] + mult_out_21[88] + mult_out_22[88])%3329) ;
                                                                                                                                       mul_add[2][89]<=((mult_out_20[89] + mult_out_21[89] + mult_out_22[89])%3329) ;
                                                                                                                                       mul_add[2][90]<=((mult_out_20[90] + mult_out_21[90] + mult_out_22[90])%3329) ;
                                                                                                                                       mul_add[2][91]<=((mult_out_20[91] + mult_out_21[91] + mult_out_22[91])%3329) ;
                                                                                                                                       mul_add[2][92]<=((mult_out_20[92] + mult_out_21[92] + mult_out_22[92])%3329) ;
                                                                                                                                       mul_add[2][93]<=((mult_out_20[93] + mult_out_21[93] + mult_out_22[93])%3329) ;
                                                                                                                                       mul_add[2][94]<=((mult_out_20[94] + mult_out_21[94] + mult_out_22[94])%3329) ;
                                                                                                                                       mul_add[2][95]<=((mult_out_20[95] + mult_out_21[95] + mult_out_22[95])%3329) ;
                                                                                                                                       mul_add[2][96]<=((mult_out_20[96] + mult_out_21[96] + mult_out_22[96])%3329) ;
                                                                                                                                       mul_add[2][97]<=((mult_out_20[97] + mult_out_21[97] + mult_out_22[97])%3329) ;
                                                                                                                                       mul_add[2][98]<=((mult_out_20[98] + mult_out_21[98] + mult_out_22[98])%3329) ;
                                                                                                                                       mul_add[2][99]<=((mult_out_20[99] + mult_out_21[99] + mult_out_22[99])%3329) ;
                                                                                                                                       mul_add[2][100]<=((mult_out_20[100] + mult_out_21[100] + mult_out_22[100])%3329) ;
                                                                                                                                       mul_add[2][101]<=((mult_out_20[101] + mult_out_21[101] + mult_out_22[101])%3329) ;
                                                                                                                                       mul_add[2][102]<=((mult_out_20[102] + mult_out_21[102] + mult_out_22[102])%3329) ;
                                                                                                                                       mul_add[2][103]<=((mult_out_20[103] + mult_out_21[103] + mult_out_22[103])%3329) ;
                                                                                                                                       mul_add[2][104]<=((mult_out_20[104] + mult_out_21[104] + mult_out_22[104])%3329) ;
                                                                                                                                       mul_add[2][105]<=((mult_out_20[105] + mult_out_21[105] + mult_out_22[105])%3329) ;
                                                                                                                                       mul_add[2][106]<=((mult_out_20[106] + mult_out_21[106] + mult_out_22[106])%3329) ;
                                                                                                                                       mul_add[2][107]<=((mult_out_20[107] + mult_out_21[107] + mult_out_22[107])%3329) ;
                                                                                                                                       mul_add[2][108]<=((mult_out_20[108] + mult_out_21[108] + mult_out_22[108])%3329) ;
                                                                                                                                       mul_add[2][109]<=((mult_out_20[109] + mult_out_21[109] + mult_out_22[109])%3329) ;
                                                                                                                                       mul_add[2][110]<=((mult_out_20[110] + mult_out_21[110] + mult_out_22[110])%3329) ;
                                                                                                                                       mul_add[2][111]<=((mult_out_20[111] + mult_out_21[111] + mult_out_22[111])%3329) ;
                                                                                                                                       mul_add[2][112]<=((mult_out_20[112] + mult_out_21[112] + mult_out_22[112])%3329) ;
                                                                                                                                       mul_add[2][113]<=((mult_out_20[113] + mult_out_21[113] + mult_out_22[113])%3329) ;
                                                                                                                                       mul_add[2][114]<=((mult_out_20[114] + mult_out_21[114] + mult_out_22[114])%3329) ;
                                                                                                                                       mul_add[2][115]<=((mult_out_20[115] + mult_out_21[115] + mult_out_22[115])%3329) ;
                                                                                                                                       mul_add[2][116]<=((mult_out_20[116] + mult_out_21[116] + mult_out_22[116])%3329) ;
                                                                                                                                       mul_add[2][117]<=((mult_out_20[117] + mult_out_21[117] + mult_out_22[117])%3329) ;
                                                                                                                                       mul_add[2][118]<=((mult_out_20[118] + mult_out_21[118] + mult_out_22[118])%3329) ;
                                                                                                                                       mul_add[2][119]<=((mult_out_20[119] + mult_out_21[119] + mult_out_22[119])%3329) ;
                                                                                                                                       mul_add[2][120]<=((mult_out_20[120] + mult_out_21[120] + mult_out_22[120])%3329) ;
                                                                                                                                       mul_add[2][121]<=((mult_out_20[121] + mult_out_21[121] + mult_out_22[121])%3329) ;
                                                                                                                                       mul_add[2][122]<=((mult_out_20[122] + mult_out_21[122] + mult_out_22[122])%3329) ;
                                                                                                                                       mul_add[2][123]<=((mult_out_20[123] + mult_out_21[123] + mult_out_22[123])%3329) ;
                                                                                                                                       mul_add[2][124]<=((mult_out_20[124] + mult_out_21[124] + mult_out_22[124])%3329) ;
                                                                                                                                       mul_add[2][125]<=((mult_out_20[125] + mult_out_21[125] + mult_out_22[125])%3329) ;
                                                                                                                                       mul_add[2][126]<=((mult_out_20[126] + mult_out_21[126] + mult_out_22[126])%3329) ;
                                                                                                                                       mul_add[2][127]<=((mult_out_20[127] + mult_out_21[127] + mult_out_22[127])%3329) ;
                                                                                                                                       mul_add[2][128]<=((mult_out_20[128] + mult_out_21[128] + mult_out_22[128])%3329) ;
                                                                                                                                       mul_add[2][129]<=((mult_out_20[129] + mult_out_21[129] + mult_out_22[129])%3329) ;
                                                                                                                                       mul_add[2][130]<=((mult_out_20[130] + mult_out_21[130] + mult_out_22[130])%3329) ;
                                                                                                                                       mul_add[2][131]<=((mult_out_20[131] + mult_out_21[131] + mult_out_22[131])%3329) ;
                                                                                                                                       mul_add[2][132]<=((mult_out_20[132] + mult_out_21[132] + mult_out_22[132])%3329) ;
                                                                                                                                       mul_add[2][133]<=((mult_out_20[133] + mult_out_21[133] + mult_out_22[133])%3329) ;
                                                                                                                                       mul_add[2][134]<=((mult_out_20[134] + mult_out_21[134] + mult_out_22[134])%3329) ;
                                                                                                                                       mul_add[2][135]<=((mult_out_20[135] + mult_out_21[135] + mult_out_22[135])%3329) ;
                                                                                                                                       mul_add[2][136]<=((mult_out_20[136] + mult_out_21[136] + mult_out_22[136])%3329) ;
                                                                                                                                       mul_add[2][137]<=((mult_out_20[137] + mult_out_21[137] + mult_out_22[137])%3329) ;
                                                                                                                                       mul_add[2][138]<=((mult_out_20[138] + mult_out_21[138] + mult_out_22[138])%3329) ;
                                                                                                                                       mul_add[2][139]<=((mult_out_20[139] + mult_out_21[139] + mult_out_22[139])%3329) ;
                                                                                                                                       mul_add[2][140]<=((mult_out_20[140] + mult_out_21[140] + mult_out_22[140])%3329) ;
                                                                                                                                       mul_add[2][141]<=((mult_out_20[141] + mult_out_21[141] + mult_out_22[141])%3329) ;
                                                                                                                                       mul_add[2][142]<=((mult_out_20[142] + mult_out_21[142] + mult_out_22[142])%3329) ;
                                                                                                                                       mul_add[2][143]<=((mult_out_20[143] + mult_out_21[143] + mult_out_22[143])%3329) ;
                                                                                                                                       mul_add[2][144]<=((mult_out_20[144] + mult_out_21[144] + mult_out_22[144])%3329) ;
                                                                                                                                       mul_add[2][145]<=((mult_out_20[145] + mult_out_21[145] + mult_out_22[145])%3329) ;
                                                                                                                                       mul_add[2][146]<=((mult_out_20[146] + mult_out_21[146] + mult_out_22[146])%3329) ;
                                                                                                                                       mul_add[2][147]<=((mult_out_20[147] + mult_out_21[147] + mult_out_22[147])%3329) ;
                                                                                                                                       mul_add[2][148]<=((mult_out_20[148] + mult_out_21[148] + mult_out_22[148])%3329) ;
                                                                                                                                       mul_add[2][149]<=((mult_out_20[149] + mult_out_21[149] + mult_out_22[149])%3329) ;
                                                                                                                                       mul_add[2][150]<=((mult_out_20[150] + mult_out_21[150] + mult_out_22[150])%3329) ;
                                                                                                                                       mul_add[2][151]<=((mult_out_20[151] + mult_out_21[151] + mult_out_22[151])%3329) ;
                                                                                                                                       mul_add[2][152]<=((mult_out_20[152] + mult_out_21[152] + mult_out_22[152])%3329) ;
                                                                                                                                       mul_add[2][153]<=((mult_out_20[153] + mult_out_21[153] + mult_out_22[153])%3329) ;
                                                                                                                                       mul_add[2][154]<=((mult_out_20[154] + mult_out_21[154] + mult_out_22[154])%3329) ;
                                                                                                                                       mul_add[2][155]<=((mult_out_20[155] + mult_out_21[155] + mult_out_22[155])%3329) ;
                                                                                                                                       mul_add[2][156]<=((mult_out_20[156] + mult_out_21[156] + mult_out_22[156])%3329) ;
                                                                                                                                       mul_add[2][157]<=((mult_out_20[157] + mult_out_21[157] + mult_out_22[157])%3329) ;
                                                                                                                                       mul_add[2][158]<=((mult_out_20[158] + mult_out_21[158] + mult_out_22[158])%3329) ;
                                                                                                                                       mul_add[2][159]<=((mult_out_20[159] + mult_out_21[159] + mult_out_22[159])%3329) ;
                                                                                                                                       mul_add[2][160]<=((mult_out_20[160] + mult_out_21[160] + mult_out_22[160])%3329) ;
                                                                                                                                       mul_add[2][161]<=((mult_out_20[161] + mult_out_21[161] + mult_out_22[161])%3329) ;
                                                                                                                                       mul_add[2][162]<=((mult_out_20[162] + mult_out_21[162] + mult_out_22[162])%3329) ;
                                                                                                                                       mul_add[2][163]<=((mult_out_20[163] + mult_out_21[163] + mult_out_22[163])%3329) ;
                                                                                                                                       mul_add[2][164]<=((mult_out_20[164] + mult_out_21[164] + mult_out_22[164])%3329) ;
                                                                                                                                       mul_add[2][165]<=((mult_out_20[165] + mult_out_21[165] + mult_out_22[165])%3329) ;
                                                                                                                                       mul_add[2][166]<=((mult_out_20[166] + mult_out_21[166] + mult_out_22[166])%3329) ;
                                                                                                                                       mul_add[2][167]<=((mult_out_20[167] + mult_out_21[167] + mult_out_22[167])%3329) ;
                                                                                                                                       mul_add[2][168]<=((mult_out_20[168] + mult_out_21[168] + mult_out_22[168])%3329) ;
                                                                                                                                       mul_add[2][169]<=((mult_out_20[169] + mult_out_21[169] + mult_out_22[169])%3329) ;
                                                                                                                                       mul_add[2][170]<=((mult_out_20[170] + mult_out_21[170] + mult_out_22[170])%3329) ;
                                                                                                                                       mul_add[2][171]<=((mult_out_20[171] + mult_out_21[171] + mult_out_22[171])%3329) ;
                                                                                                                                       mul_add[2][172]<=((mult_out_20[172] + mult_out_21[172] + mult_out_22[172])%3329) ;
                                                                                                                                       mul_add[2][173]<=((mult_out_20[173] + mult_out_21[173] + mult_out_22[173])%3329) ;
                                                                                                                                       mul_add[2][174]<=((mult_out_20[174] + mult_out_21[174] + mult_out_22[174])%3329) ;
                                                                                                                                       mul_add[2][175]<=((mult_out_20[175] + mult_out_21[175] + mult_out_22[175])%3329) ;
                                                                                                                                       mul_add[2][176]<=((mult_out_20[176] + mult_out_21[176] + mult_out_22[176])%3329) ;
                                                                                                                                       mul_add[2][177]<=((mult_out_20[177] + mult_out_21[177] + mult_out_22[177])%3329) ;
                                                                                                                                       mul_add[2][178]<=((mult_out_20[178] + mult_out_21[178] + mult_out_22[178])%3329) ;
                                                                                                                                       mul_add[2][179]<=((mult_out_20[179] + mult_out_21[179] + mult_out_22[179])%3329) ;
                                                                                                                                       mul_add[2][180]<=((mult_out_20[180] + mult_out_21[180] + mult_out_22[180])%3329) ;
                                                                                                                                       mul_add[2][181]<=((mult_out_20[181] + mult_out_21[181] + mult_out_22[181])%3329) ;
                                                                                                                                       mul_add[2][182]<=((mult_out_20[182] + mult_out_21[182] + mult_out_22[182])%3329) ;
                                                                                                                                       mul_add[2][183]<=((mult_out_20[183] + mult_out_21[183] + mult_out_22[183])%3329) ;
                                                                                                                                       mul_add[2][184]<=((mult_out_20[184] + mult_out_21[184] + mult_out_22[184])%3329) ;
                                                                                                                                       mul_add[2][185]<=((mult_out_20[185] + mult_out_21[185] + mult_out_22[185])%3329) ;
                                                                                                                                       mul_add[2][186]<=((mult_out_20[186] + mult_out_21[186] + mult_out_22[186])%3329) ;
                                                                                                                                       mul_add[2][187]<=((mult_out_20[187] + mult_out_21[187] + mult_out_22[187])%3329) ;
                                                                                                                                       mul_add[2][188]<=((mult_out_20[188] + mult_out_21[188] + mult_out_22[188])%3329) ;
                                                                                                                                       mul_add[2][189]<=((mult_out_20[189] + mult_out_21[189] + mult_out_22[189])%3329) ;
                                                                                                                                       mul_add[2][190]<=((mult_out_20[190] + mult_out_21[190] + mult_out_22[190])%3329) ;
                                                                                                                                       mul_add[2][191]<=((mult_out_20[191] + mult_out_21[191] + mult_out_22[191])%3329) ;
                                                                                                                                       mul_add[2][192]<=((mult_out_20[192] + mult_out_21[192] + mult_out_22[192])%3329) ;
                                                                                                                                       mul_add[2][193]<=((mult_out_20[193] + mult_out_21[193] + mult_out_22[193])%3329) ;
                                                                                                                                       mul_add[2][194]<=((mult_out_20[194] + mult_out_21[194] + mult_out_22[194])%3329) ;
                                                                                                                                       mul_add[2][195]<=((mult_out_20[195] + mult_out_21[195] + mult_out_22[195])%3329) ;
                                                                                                                                       mul_add[2][196]<=((mult_out_20[196] + mult_out_21[196] + mult_out_22[196])%3329) ;
                                                                                                                                       mul_add[2][197]<=((mult_out_20[197] + mult_out_21[197] + mult_out_22[197])%3329) ;
                                                                                                                                       mul_add[2][198]<=((mult_out_20[198] + mult_out_21[198] + mult_out_22[198])%3329) ;
                                                                                                                                       mul_add[2][199]<=((mult_out_20[199] + mult_out_21[199] + mult_out_22[199])%3329) ;
                                                                                                                                       mul_add[2][200]<=((mult_out_20[200] + mult_out_21[200] + mult_out_22[200])%3329) ;
                                                                                                                                       mul_add[2][201]<=((mult_out_20[201] + mult_out_21[201] + mult_out_22[201])%3329) ;
                                                                                                                                       mul_add[2][202]<=((mult_out_20[202] + mult_out_21[202] + mult_out_22[202])%3329) ;
                                                                                                                                       mul_add[2][203]<=((mult_out_20[203] + mult_out_21[203] + mult_out_22[203])%3329) ;
                                                                                                                                       mul_add[2][204]<=((mult_out_20[204] + mult_out_21[204] + mult_out_22[204])%3329) ;
                                                                                                                                       mul_add[2][205]<=((mult_out_20[205] + mult_out_21[205] + mult_out_22[205])%3329) ;
                                                                                                                                       mul_add[2][206]<=((mult_out_20[206] + mult_out_21[206] + mult_out_22[206])%3329) ;
                                                                                                                                       mul_add[2][207]<=((mult_out_20[207] + mult_out_21[207] + mult_out_22[207])%3329) ;
                                                                                                                                       mul_add[2][208]<=((mult_out_20[208] + mult_out_21[208] + mult_out_22[208])%3329) ;
                                                                                                                                       mul_add[2][209]<=((mult_out_20[209] + mult_out_21[209] + mult_out_22[209])%3329) ;
                                                                                                                                       mul_add[2][210]<=((mult_out_20[210] + mult_out_21[210] + mult_out_22[210])%3329) ;
                                                                                                                                       mul_add[2][211]<=((mult_out_20[211] + mult_out_21[211] + mult_out_22[211])%3329) ;
                                                                                                                                       mul_add[2][212]<=((mult_out_20[212] + mult_out_21[212] + mult_out_22[212])%3329) ;
                                                                                                                                       mul_add[2][213]<=((mult_out_20[213] + mult_out_21[213] + mult_out_22[213])%3329) ;
                                                                                                                                       mul_add[2][214]<=((mult_out_20[214] + mult_out_21[214] + mult_out_22[214])%3329) ;
                                                                                                                                       mul_add[2][215]<=((mult_out_20[215] + mult_out_21[215] + mult_out_22[215])%3329) ;
                                                                                                                                       mul_add[2][216]<=((mult_out_20[216] + mult_out_21[216] + mult_out_22[216])%3329) ;
                                                                                                                                       mul_add[2][217]<=((mult_out_20[217] + mult_out_21[217] + mult_out_22[217])%3329) ;
                                                                                                                                       mul_add[2][218]<=((mult_out_20[218] + mult_out_21[218] + mult_out_22[218])%3329) ;
                                                                                                                                       mul_add[2][219]<=((mult_out_20[219] + mult_out_21[219] + mult_out_22[219])%3329) ;
                                                                                                                                       mul_add[2][220]<=((mult_out_20[220] + mult_out_21[220] + mult_out_22[220])%3329) ;
                                                                                                                                       mul_add[2][221]<=((mult_out_20[221] + mult_out_21[221] + mult_out_22[221])%3329) ;
                                                                                                                                       mul_add[2][222]<=((mult_out_20[222] + mult_out_21[222] + mult_out_22[222])%3329) ;
                                                                                                                                       mul_add[2][223]<=((mult_out_20[223] + mult_out_21[223] + mult_out_22[223])%3329) ;
                                                                                                                                       mul_add[2][224]<=((mult_out_20[224] + mult_out_21[224] + mult_out_22[224])%3329) ;
                                                                                                                                       mul_add[2][225]<=((mult_out_20[225] + mult_out_21[225] + mult_out_22[225])%3329) ;
                                                                                                                                       mul_add[2][226]<=((mult_out_20[226] + mult_out_21[226] + mult_out_22[226])%3329) ;
                                                                                                                                       mul_add[2][227]<=((mult_out_20[227] + mult_out_21[227] + mult_out_22[227])%3329) ;
                                                                                                                                       mul_add[2][228]<=((mult_out_20[228] + mult_out_21[228] + mult_out_22[228])%3329) ;
                                                                                                                                       mul_add[2][229]<=((mult_out_20[229] + mult_out_21[229] + mult_out_22[229])%3329) ;
                                                                                                                                       mul_add[2][230]<=((mult_out_20[230] + mult_out_21[230] + mult_out_22[230])%3329) ;
                                                                                                                                       mul_add[2][231]<=((mult_out_20[231] + mult_out_21[231] + mult_out_22[231])%3329) ;
                                                                                                                                       mul_add[2][232]<=((mult_out_20[232] + mult_out_21[232] + mult_out_22[232])%3329) ;
                                                                                                                                       mul_add[2][233]<=((mult_out_20[233] + mult_out_21[233] + mult_out_22[233])%3329) ;
                                                                                                                                       mul_add[2][234]<=((mult_out_20[234] + mult_out_21[234] + mult_out_22[234])%3329) ;
                                                                                                                                       mul_add[2][235]<=((mult_out_20[235] + mult_out_21[235] + mult_out_22[235])%3329) ;
                                                                                                                                       mul_add[2][236]<=((mult_out_20[236] + mult_out_21[236] + mult_out_22[236])%3329) ;
                                                                                                                                       mul_add[2][237]<=((mult_out_20[237] + mult_out_21[237] + mult_out_22[237])%3329) ;
                                                                                                                                       mul_add[2][238]<=((mult_out_20[238] + mult_out_21[238] + mult_out_22[238])%3329) ;
                                                                                                                                       mul_add[2][239]<=((mult_out_20[239] + mult_out_21[239] + mult_out_22[239])%3329) ;
                                                                                                                                       mul_add[2][240]<=((mult_out_20[240] + mult_out_21[240] + mult_out_22[240])%3329) ;
                                                                                                                                       mul_add[2][241]<=((mult_out_20[241] + mult_out_21[241] + mult_out_22[241])%3329) ;
                                                                                                                                       mul_add[2][242]<=((mult_out_20[242] + mult_out_21[242] + mult_out_22[242])%3329) ;
                                                                                                                                       mul_add[2][243]<=((mult_out_20[243] + mult_out_21[243] + mult_out_22[243])%3329) ;
                                                                                                                                       mul_add[2][244]<=((mult_out_20[244] + mult_out_21[244] + mult_out_22[244])%3329) ;
                                                                                                                                       mul_add[2][245]<=((mult_out_20[245] + mult_out_21[245] + mult_out_22[245])%3329) ;
                                                                                                                                       mul_add[2][246]<=((mult_out_20[246] + mult_out_21[246] + mult_out_22[246])%3329) ;
                                                                                                                                       mul_add[2][247]<=((mult_out_20[247] + mult_out_21[247] + mult_out_22[247])%3329) ;
                                                                                                                                       mul_add[2][248]<=((mult_out_20[248] + mult_out_21[248] + mult_out_22[248])%3329) ;
                                                                                                                                       mul_add[2][249]<=((mult_out_20[249] + mult_out_21[249] + mult_out_22[249])%3329) ;
                                                                                                                                       mul_add[2][250]<=((mult_out_20[250] + mult_out_21[250] + mult_out_22[250])%3329) ;
                                                                                                                                       mul_add[2][251]<=((mult_out_20[251] + mult_out_21[251] + mult_out_22[251])%3329) ;
                                                                                                                                       mul_add[2][252]<=((mult_out_20[252] + mult_out_21[252] + mult_out_22[252])%3329) ;
                                                                                                                                       mul_add[2][253]<=((mult_out_20[253] + mult_out_21[253] + mult_out_22[253])%3329) ;
                                                                                                                                       mul_add[2][254]<=((mult_out_20[254] + mult_out_21[254] + mult_out_22[254])%3329) ;
                                                                                                                                       mul_add[2][255]<=((mult_out_20[255] + mult_out_21[255] + mult_out_22[255])%3329) ;
                                                                                                                                                                                                             
                                                                                                                                                           if (done9_mul && done10_mul && done11_mul) begin
                                                                                                                                                                  mul_add_t[0][0] <= (mult_out_1[0] + mult_out_2[0] + mult_out_3[0]) % 3329;
                                                                                                                                                                  mul_add_t[0][1] <= (mult_out_1[1] + mult_out_2[1] + mult_out_3[1]) % 3329;
                                                                                                                                                                  mul_add_t[0][2] <= (mult_out_1[2] + mult_out_2[2] + mult_out_3[2]) % 3329;
                                                                                                                                                                  mul_add_t[0][3] <= (mult_out_1[3] + mult_out_2[3] + mult_out_3[3]) % 3329;
                                                                                                                                                                  mul_add_t[0][4] <= (mult_out_1[4] + mult_out_2[4] + mult_out_3[4]) % 3329;
                                                                                                                                                                  mul_add_t[0][5] <= (mult_out_1[5] + mult_out_2[5] + mult_out_3[5]) % 3329;
                                                                                                                                                                  mul_add_t[0][6] <= (mult_out_1[6] + mult_out_2[6] + mult_out_3[6]) % 3329;
                                                                                                                                                                  mul_add_t[0][7] <= (mult_out_1[7] + mult_out_2[7] + mult_out_3[7]) % 3329;
                                                                                                                                                                  mul_add_t[0][8] <= (mult_out_1[8] + mult_out_2[8] + mult_out_3[8]) % 3329;
                                                                                                                                                                  mul_add_t[0][9] <= (mult_out_1[9] + mult_out_2[9] + mult_out_3[9]) % 3329;
                                                                                                                                                                  mul_add_t[0][10] <= (mult_out_1[10] + mult_out_2[10] + mult_out_3[10]) % 3329;
                                                                                                                                                                  mul_add_t[0][11] <= (mult_out_1[11] + mult_out_2[11] + mult_out_3[11]) % 3329;
                                                                                                                                                                  mul_add_t[0][12] <= (mult_out_1[12] + mult_out_2[12] + mult_out_3[12]) % 3329;
                                                                                                                                                                  mul_add_t[0][13] <= (mult_out_1[13] + mult_out_2[13] + mult_out_3[13]) % 3329;
                                                                                                                                                                  mul_add_t[0][14] <= (mult_out_1[14] + mult_out_2[14] + mult_out_3[14]) % 3329;
                                                                                                                                                                  mul_add_t[0][15] <= (mult_out_1[15] + mult_out_2[15] + mult_out_3[15]) % 3329;
                                                                                                                                                                  mul_add_t[0][16] <= (mult_out_1[16] + mult_out_2[16] + mult_out_3[16]) % 3329;
                                                                                                                                                                  mul_add_t[0][17] <= (mult_out_1[17] + mult_out_2[17] + mult_out_3[17]) % 3329;
                                                                                                                                                                  mul_add_t[0][18] <= (mult_out_1[18] + mult_out_2[18] + mult_out_3[18]) % 3329;
                                                                                                                                                                  mul_add_t[0][19] <= (mult_out_1[19] + mult_out_2[19] + mult_out_3[19]) % 3329;
                                                                                                                                                                  mul_add_t[0][20] <= (mult_out_1[20] + mult_out_2[20] + mult_out_3[20]) % 3329;
                                                                                                                                                                  mul_add_t[0][21] <= (mult_out_1[21] + mult_out_2[21] + mult_out_3[21]) % 3329;
                                                                                                                                                                  mul_add_t[0][22] <= (mult_out_1[22] + mult_out_2[22] + mult_out_3[22]) % 3329;
                                                                                                                                                                  mul_add_t[0][23] <= (mult_out_1[23] + mult_out_2[23] + mult_out_3[23]) % 3329;
                                                                                                                                                                  mul_add_t[0][24] <= (mult_out_1[24] + mult_out_2[24] + mult_out_3[24]) % 3329;
                                                                                                                                                                  mul_add_t[0][25] <= (mult_out_1[25] + mult_out_2[25] + mult_out_3[25]) % 3329;
                                                                                                                                                                  mul_add_t[0][26] <= (mult_out_1[26] + mult_out_2[26] + mult_out_3[26]) % 3329;
                                                                                                                                                                  mul_add_t[0][27] <= (mult_out_1[27] + mult_out_2[27] + mult_out_3[27]) % 3329;
                                                                                                                                                                  mul_add_t[0][28] <= (mult_out_1[28] + mult_out_2[28] + mult_out_3[28]) % 3329;
                                                                                                                                                                  mul_add_t[0][29] <= (mult_out_1[29] + mult_out_2[29] + mult_out_3[29]) % 3329;
                                                                                                                                                                  mul_add_t[0][30] <= (mult_out_1[30] + mult_out_2[30] + mult_out_3[30]) % 3329;
                                                                                                                                                                  mul_add_t[0][31] <= (mult_out_1[31] + mult_out_2[31] + mult_out_3[31]) % 3329;
                                                                                                                                                                  mul_add_t[0][32] <= (mult_out_1[32] + mult_out_2[32] + mult_out_3[32]) % 3329;
                                                                                                                                                                  mul_add_t[0][33] <= (mult_out_1[33] + mult_out_2[33] + mult_out_3[33]) % 3329;
                                                                                                                                                                  mul_add_t[0][34] <= (mult_out_1[34] + mult_out_2[34] + mult_out_3[34]) % 3329;
                                                                                                                                                                  mul_add_t[0][35] <= (mult_out_1[35] + mult_out_2[35] + mult_out_3[35]) % 3329;
                                                                                                                                                                  mul_add_t[0][36] <= (mult_out_1[36] + mult_out_2[36] + mult_out_3[36]) % 3329;
                                                                                                                                                                  mul_add_t[0][37] <= (mult_out_1[37] + mult_out_2[37] + mult_out_3[37]) % 3329;
                                                                                                                                                                  mul_add_t[0][38] <= (mult_out_1[38] + mult_out_2[38] + mult_out_3[38]) % 3329;
                                                                                                                                                                  mul_add_t[0][39] <= (mult_out_1[39] + mult_out_2[39] + mult_out_3[39]) % 3329;
                                                                                                                                                                  mul_add_t[0][40] <= (mult_out_1[40] + mult_out_2[40] + mult_out_3[40]) % 3329;
                                                                                                                                                                  mul_add_t[0][41] <= (mult_out_1[41] + mult_out_2[41] + mult_out_3[41]) % 3329;
                                                                                                                                                                  mul_add_t[0][42] <= (mult_out_1[42] + mult_out_2[42] + mult_out_3[42]) % 3329;
                                                                                                                                                                  mul_add_t[0][43] <= (mult_out_1[43] + mult_out_2[43] + mult_out_3[43]) % 3329;
                                                                                                                                                                  mul_add_t[0][44] <= (mult_out_1[44] + mult_out_2[44] + mult_out_3[44]) % 3329;
                                                                                                                                                                  mul_add_t[0][45] <= (mult_out_1[45] + mult_out_2[45] + mult_out_3[45]) % 3329;
                                                                                                                                                                  mul_add_t[0][46] <= (mult_out_1[46] + mult_out_2[46] + mult_out_3[46]) % 3329;
                                                                                                                                                                  mul_add_t[0][47] <= (mult_out_1[47] + mult_out_2[47] + mult_out_3[47]) % 3329;
                                                                                                                                                                  mul_add_t[0][48] <= (mult_out_1[48] + mult_out_2[48] + mult_out_3[48]) % 3329;
                                                                                                                                                                  mul_add_t[0][49] <= (mult_out_1[49] + mult_out_2[49] + mult_out_3[49]) % 3329;
                                                                                                                                                                  mul_add_t[0][50] <= (mult_out_1[50] + mult_out_2[50] + mult_out_3[50]) % 3329;
                                                                                                                                                                  mul_add_t[0][51] <= (mult_out_1[51] + mult_out_2[51] + mult_out_3[51]) % 3329;
                                                                                                                                                                  mul_add_t[0][52] <= (mult_out_1[52] + mult_out_2[52] + mult_out_3[52]) % 3329;
                                                                                                                                                                  mul_add_t[0][53] <= (mult_out_1[53] + mult_out_2[53] + mult_out_3[53]) % 3329;
                                                                                                                                                                  mul_add_t[0][54] <= (mult_out_1[54] + mult_out_2[54] + mult_out_3[54]) % 3329;
                                                                                                                                                                  mul_add_t[0][55] <= (mult_out_1[55] + mult_out_2[55] + mult_out_3[55]) % 3329;
                                                                                                                                                                  mul_add_t[0][56] <= (mult_out_1[56] + mult_out_2[56] + mult_out_3[56]) % 3329;
                                                                                                                                                                  mul_add_t[0][57] <= (mult_out_1[57] + mult_out_2[57] + mult_out_3[57]) % 3329;
                                                                                                                                                                  mul_add_t[0][58] <= (mult_out_1[58] + mult_out_2[58] + mult_out_3[58]) % 3329;
                                                                                                                                                                  mul_add_t[0][59] <= (mult_out_1[59] + mult_out_2[59] + mult_out_3[59]) % 3329;
                                                                                                                                                                  mul_add_t[0][60] <= (mult_out_1[60] + mult_out_2[60] + mult_out_3[60]) % 3329;
                                                                                                                                                                  mul_add_t[0][61] <= (mult_out_1[61] + mult_out_2[61] + mult_out_3[61]) % 3329;
                                                                                                                                                                  mul_add_t[0][62] <= (mult_out_1[62] + mult_out_2[62] + mult_out_3[62]) % 3329;
                                                                                                                                                                  mul_add_t[0][63] <= (mult_out_1[63] + mult_out_2[63] + mult_out_3[63]) % 3329;
                                                                                                                                                                  mul_add_t[0][64] <= (mult_out_1[64] + mult_out_2[64] + mult_out_3[64]) % 3329;
                                                                                                                                                                  mul_add_t[0][65] <= (mult_out_1[65] + mult_out_2[65] + mult_out_3[65]) % 3329;
                                                                                                                                                                  mul_add_t[0][66] <= (mult_out_1[66] + mult_out_2[66] + mult_out_3[66]) % 3329;
                                                                                                                                                                  mul_add_t[0][67] <= (mult_out_1[67] + mult_out_2[67] + mult_out_3[67]) % 3329;
                                                                                                                                                                  mul_add_t[0][68] <= (mult_out_1[68] + mult_out_2[68] + mult_out_3[68]) % 3329;
                                                                                                                                                                  mul_add_t[0][69] <= (mult_out_1[69] + mult_out_2[69] + mult_out_3[69]) % 3329;
                                                                                                                                                                  mul_add_t[0][70] <= (mult_out_1[70] + mult_out_2[70] + mult_out_3[70]) % 3329;
                                                                                                                                                                  mul_add_t[0][71] <= (mult_out_1[71] + mult_out_2[71] + mult_out_3[71]) % 3329;
                                                                                                                                                                  mul_add_t[0][72] <= (mult_out_1[72] + mult_out_2[72] + mult_out_3[72]) % 3329;
                                                                                                                                                                  mul_add_t[0][73] <= (mult_out_1[73] + mult_out_2[73] + mult_out_3[73]) % 3329;
                                                                                                                                                                  mul_add_t[0][74] <= (mult_out_1[74] + mult_out_2[74] + mult_out_3[74]) % 3329;
                                                                                                                                                                  mul_add_t[0][75] <= (mult_out_1[75] + mult_out_2[75] + mult_out_3[75]) % 3329;
                                                                                                                                                                  mul_add_t[0][76] <= (mult_out_1[76] + mult_out_2[76] + mult_out_3[76]) % 3329;
                                                                                                                                                                  mul_add_t[0][77] <= (mult_out_1[77] + mult_out_2[77] + mult_out_3[77]) % 3329;
                                                                                                                                                                  mul_add_t[0][78] <= (mult_out_1[78] + mult_out_2[78] + mult_out_3[78]) % 3329;
                                                                                                                                                                  mul_add_t[0][79] <= (mult_out_1[79] + mult_out_2[79] + mult_out_3[79]) % 3329;
                                                                                                                                                                  mul_add_t[0][80] <= (mult_out_1[80] + mult_out_2[80] + mult_out_3[80]) % 3329;
                                                                                                                                                                  mul_add_t[0][81] <= (mult_out_1[81] + mult_out_2[81] + mult_out_3[81]) % 3329;
                                                                                                                                                                  mul_add_t[0][82] <= (mult_out_1[82] + mult_out_2[82] + mult_out_3[82]) % 3329;
                                                                                                                                                                  mul_add_t[0][83] <= (mult_out_1[83] + mult_out_2[83] + mult_out_3[83]) % 3329;
                                                                                                                                                                  mul_add_t[0][84] <= (mult_out_1[84] + mult_out_2[84] + mult_out_3[84]) % 3329;
                                                                                                                                                                  mul_add_t[0][85] <= (mult_out_1[85] + mult_out_2[85] + mult_out_3[85]) % 3329;
                                                                                                                                                                  mul_add_t[0][86] <= (mult_out_1[86] + mult_out_2[86] + mult_out_3[86]) % 3329;
                                                                                                                                                                  mul_add_t[0][87] <= (mult_out_1[87] + mult_out_2[87] + mult_out_3[87]) % 3329;
                                                                                                                                                                  mul_add_t[0][88] <= (mult_out_1[88] + mult_out_2[88] + mult_out_3[88]) % 3329;
                                                                                                                                                                  mul_add_t[0][89] <= (mult_out_1[89] + mult_out_2[89] + mult_out_3[89]) % 3329;
                                                                                                                                                                  mul_add_t[0][90] <= (mult_out_1[90] + mult_out_2[90] + mult_out_3[90]) % 3329;
                                                                                                                                                                  mul_add_t[0][91] <= (mult_out_1[91] + mult_out_2[91] + mult_out_3[91]) % 3329;
                                                                                                                                                                  mul_add_t[0][92] <= (mult_out_1[92] + mult_out_2[92] + mult_out_3[92]) % 3329;
                                                                                                                                                                  mul_add_t[0][93] <= (mult_out_1[93] + mult_out_2[93] + mult_out_3[93]) % 3329;
                                                                                                                                                                  mul_add_t[0][94] <= (mult_out_1[94] + mult_out_2[94] + mult_out_3[94]) % 3329;
                                                                                                                                                                  mul_add_t[0][95] <= (mult_out_1[95] + mult_out_2[95] + mult_out_3[95]) % 3329;
                                                                                                                                                                  mul_add_t[0][96] <= (mult_out_1[96] + mult_out_2[96] + mult_out_3[96]) % 3329;
                                                                                                                                                                  mul_add_t[0][97] <= (mult_out_1[97] + mult_out_2[97] + mult_out_3[97]) % 3329;
                                                                                                                                                                  mul_add_t[0][98] <= (mult_out_1[98] + mult_out_2[98] + mult_out_3[98]) % 3329;
                                                                                                                                                                  mul_add_t[0][99] <= (mult_out_1[99] + mult_out_2[99] + mult_out_3[99]) % 3329;
                                                                                                                                                                  mul_add_t[0][100] <= (mult_out_1[100] + mult_out_2[100] + mult_out_3[100]) % 3329;
                                                                                                                                                                  mul_add_t[0][101] <= (mult_out_1[101] + mult_out_2[101] + mult_out_3[101]) % 3329;
                                                                                                                                                                  mul_add_t[0][102] <= (mult_out_1[102] + mult_out_2[102] + mult_out_3[102]) % 3329;
                                                                                                                                                                  mul_add_t[0][103] <= (mult_out_1[103] + mult_out_2[103] + mult_out_3[103]) % 3329;
                                                                                                                                                                  mul_add_t[0][104] <= (mult_out_1[104] + mult_out_2[104] + mult_out_3[104]) % 3329;
                                                                                                                                                                  mul_add_t[0][105] <= (mult_out_1[105] + mult_out_2[105] + mult_out_3[105]) % 3329;
                                                                                                                                                                  mul_add_t[0][106] <= (mult_out_1[106] + mult_out_2[106] + mult_out_3[106]) % 3329;
                                                                                                                                                                  mul_add_t[0][107] <= (mult_out_1[107] + mult_out_2[107] + mult_out_3[107]) % 3329;
                                                                                                                                                                  mul_add_t[0][108] <= (mult_out_1[108] + mult_out_2[108] + mult_out_3[108]) % 3329;
                                                                                                                                                                  mul_add_t[0][109] <= (mult_out_1[109] + mult_out_2[109] + mult_out_3[109]) % 3329;
                                                                                                                                                                  mul_add_t[0][110] <= (mult_out_1[110] + mult_out_2[110] + mult_out_3[110]) % 3329;
                                                                                                                                                                  mul_add_t[0][111] <= (mult_out_1[111] + mult_out_2[111] + mult_out_3[111]) % 3329;
                                                                                                                                                                  mul_add_t[0][112] <= (mult_out_1[112] + mult_out_2[112] + mult_out_3[112]) % 3329;
                                                                                                                                                                  mul_add_t[0][113] <= (mult_out_1[113] + mult_out_2[113] + mult_out_3[113]) % 3329;
                                                                                                                                                                  mul_add_t[0][114] <= (mult_out_1[114] + mult_out_2[114] + mult_out_3[114]) % 3329;
                                                                                                                                                                  mul_add_t[0][115] <= (mult_out_1[115] + mult_out_2[115] + mult_out_3[115]) % 3329;
                                                                                                                                                                  mul_add_t[0][116] <= (mult_out_1[116] + mult_out_2[116] + mult_out_3[116]) % 3329;
                                                                                                                                                                  mul_add_t[0][117] <= (mult_out_1[117] + mult_out_2[117] + mult_out_3[117]) % 3329;
                                                                                                                                                                  mul_add_t[0][118] <= (mult_out_1[118] + mult_out_2[118] + mult_out_3[118]) % 3329;
                                                                                                                                                                  mul_add_t[0][119] <= (mult_out_1[119] + mult_out_2[119] + mult_out_3[119]) % 3329;
                                                                                                                                                                  mul_add_t[0][120] <= (mult_out_1[120] + mult_out_2[120] + mult_out_3[120]) % 3329;
                                                                                                                                                                  mul_add_t[0][121] <= (mult_out_1[121] + mult_out_2[121] + mult_out_3[121]) % 3329;
                                                                                                                                                                  mul_add_t[0][122] <= (mult_out_1[122] + mult_out_2[122] + mult_out_3[122]) % 3329;
                                                                                                                                                                  mul_add_t[0][123] <= (mult_out_1[123] + mult_out_2[123] + mult_out_3[123]) % 3329;
                                                                                                                                                                  mul_add_t[0][124] <= (mult_out_1[124] + mult_out_2[124] + mult_out_3[124]) % 3329;
                                                                                                                                                                  mul_add_t[0][125] <= (mult_out_1[125] + mult_out_2[125] + mult_out_3[125]) % 3329;
                                                                                                                                                                  mul_add_t[0][126] <= (mult_out_1[126] + mult_out_2[126] + mult_out_3[126]) % 3329;
                                                                                                                                                                  mul_add_t[0][127] <= (mult_out_1[127] + mult_out_2[127] + mult_out_3[127]) % 3329;
                                                                                                                                                                  mul_add_t[0][128] <= (mult_out_1[128] + mult_out_2[128] + mult_out_3[128]) % 3329;
                                                                                                                                                                  mul_add_t[0][129] <= (mult_out_1[129] + mult_out_2[129] + mult_out_3[129]) % 3329;
                                                                                                                                                                  mul_add_t[0][130] <= (mult_out_1[130] + mult_out_2[130] + mult_out_3[130]) % 3329;
                                                                                                                                                                  mul_add_t[0][131] <= (mult_out_1[131] + mult_out_2[131] + mult_out_3[131]) % 3329;
                                                                                                                                                                  mul_add_t[0][132] <= (mult_out_1[132] + mult_out_2[132] + mult_out_3[132]) % 3329;
                                                                                                                                                                  mul_add_t[0][133] <= (mult_out_1[133] + mult_out_2[133] + mult_out_3[133]) % 3329;
                                                                                                                                                                  mul_add_t[0][134] <= (mult_out_1[134] + mult_out_2[134] + mult_out_3[134]) % 3329;
                                                                                                                                                                  mul_add_t[0][135] <= (mult_out_1[135] + mult_out_2[135] + mult_out_3[135]) % 3329;
                                                                                                                                                                  mul_add_t[0][136] <= (mult_out_1[136] + mult_out_2[136] + mult_out_3[136]) % 3329;
                                                                                                                                                                  mul_add_t[0][137] <= (mult_out_1[137] + mult_out_2[137] + mult_out_3[137]) % 3329;
                                                                                                                                                                  mul_add_t[0][138] <= (mult_out_1[138] + mult_out_2[138] + mult_out_3[138]) % 3329;
                                                                                                                                                                  mul_add_t[0][139] <= (mult_out_1[139] + mult_out_2[139] + mult_out_3[139]) % 3329;
                                                                                                                                                                  mul_add_t[0][140] <= (mult_out_1[140] + mult_out_2[140] + mult_out_3[140]) % 3329;
                                                                                                                                                                  mul_add_t[0][141] <= (mult_out_1[141] + mult_out_2[141] + mult_out_3[141]) % 3329;
                                                                                                                                                                  mul_add_t[0][142] <= (mult_out_1[142] + mult_out_2[142] + mult_out_3[142]) % 3329;
                                                                                                                                                                  mul_add_t[0][143] <= (mult_out_1[143] + mult_out_2[143] + mult_out_3[143]) % 3329;
                                                                                                                                                                  mul_add_t[0][144] <= (mult_out_1[144] + mult_out_2[144] + mult_out_3[144]) % 3329;
                                                                                                                                                                  mul_add_t[0][145] <= (mult_out_1[145] + mult_out_2[145] + mult_out_3[145]) % 3329;
                                                                                                                                                                  mul_add_t[0][146] <= (mult_out_1[146] + mult_out_2[146] + mult_out_3[146]) % 3329;
                                                                                                                                                                  mul_add_t[0][147] <= (mult_out_1[147] + mult_out_2[147] + mult_out_3[147]) % 3329;
                                                                                                                                                                  mul_add_t[0][148] <= (mult_out_1[148] + mult_out_2[148] + mult_out_3[148]) % 3329;
                                                                                                                                                                  mul_add_t[0][149] <= (mult_out_1[149] + mult_out_2[149] + mult_out_3[149]) % 3329;
                                                                                                                                                                  mul_add_t[0][150] <= (mult_out_1[150] + mult_out_2[150] + mult_out_3[150]) % 3329;
                                                                                                                                                                  mul_add_t[0][151] <= (mult_out_1[151] + mult_out_2[151] + mult_out_3[151]) % 3329;
                                                                                                                                                                  mul_add_t[0][152] <= (mult_out_1[152] + mult_out_2[152] + mult_out_3[152]) % 3329;
                                                                                                                                                                  mul_add_t[0][153] <= (mult_out_1[153] + mult_out_2[153] + mult_out_3[153]) % 3329;
                                                                                                                                                                  mul_add_t[0][154] <= (mult_out_1[154] + mult_out_2[154] + mult_out_3[154]) % 3329;
                                                                                                                                                                  mul_add_t[0][155] <= (mult_out_1[155] + mult_out_2[155] + mult_out_3[155]) % 3329;
                                                                                                                                                                  mul_add_t[0][156] <= (mult_out_1[156] + mult_out_2[156] + mult_out_3[156]) % 3329;
                                                                                                                                                                  mul_add_t[0][157] <= (mult_out_1[157] + mult_out_2[157] + mult_out_3[157]) % 3329;
                                                                                                                                                                  mul_add_t[0][158] <= (mult_out_1[158] + mult_out_2[158] + mult_out_3[158]) % 3329;
                                                                                                                                                                  mul_add_t[0][159] <= (mult_out_1[159] + mult_out_2[159] + mult_out_3[159]) % 3329;
                                                                                                                                                                  mul_add_t[0][160] <= (mult_out_1[160] + mult_out_2[160] + mult_out_3[160]) % 3329;
                                                                                                                                                                  mul_add_t[0][161] <= (mult_out_1[161] + mult_out_2[161] + mult_out_3[161]) % 3329;
                                                                                                                                                                  mul_add_t[0][162] <= (mult_out_1[162] + mult_out_2[162] + mult_out_3[162]) % 3329;
                                                                                                                                                                  mul_add_t[0][163] <= (mult_out_1[163] + mult_out_2[163] + mult_out_3[163]) % 3329;
                                                                                                                                                                  mul_add_t[0][164] <= (mult_out_1[164] + mult_out_2[164] + mult_out_3[164]) % 3329;
                                                                                                                                                                  mul_add_t[0][165] <= (mult_out_1[165] + mult_out_2[165] + mult_out_3[165]) % 3329;
                                                                                                                                                                  mul_add_t[0][166] <= (mult_out_1[166] + mult_out_2[166] + mult_out_3[166]) % 3329;
                                                                                                                                                                  mul_add_t[0][167] <= (mult_out_1[167] + mult_out_2[167] + mult_out_3[167]) % 3329;
                                                                                                                                                                  mul_add_t[0][168] <= (mult_out_1[168] + mult_out_2[168] + mult_out_3[168]) % 3329;
                                                                                                                                                                  mul_add_t[0][169] <= (mult_out_1[169] + mult_out_2[169] + mult_out_3[169]) % 3329;
                                                                                                                                                                  mul_add_t[0][170] <= (mult_out_1[170] + mult_out_2[170] + mult_out_3[170]) % 3329;
                                                                                                                                                                  mul_add_t[0][171] <= (mult_out_1[171] + mult_out_2[171] + mult_out_3[171]) % 3329;
                                                                                                                                                                  mul_add_t[0][172] <= (mult_out_1[172] + mult_out_2[172] + mult_out_3[172]) % 3329;
                                                                                                                                                                  mul_add_t[0][173] <= (mult_out_1[173] + mult_out_2[173] + mult_out_3[173]) % 3329;
                                                                                                                                                                  mul_add_t[0][174] <= (mult_out_1[174] + mult_out_2[174] + mult_out_3[174]) % 3329;
                                                                                                                                                                  mul_add_t[0][175] <= (mult_out_1[175] + mult_out_2[175] + mult_out_3[175]) % 3329;
                                                                                                                                                                  mul_add_t[0][176] <= (mult_out_1[176] + mult_out_2[176] + mult_out_3[176]) % 3329;
                                                                                                                                                                  mul_add_t[0][177] <= (mult_out_1[177] + mult_out_2[177] + mult_out_3[177]) % 3329;
                                                                                                                                                                  mul_add_t[0][178] <= (mult_out_1[178] + mult_out_2[178] + mult_out_3[178]) % 3329;
                                                                                                                                                                  mul_add_t[0][179] <= (mult_out_1[179] + mult_out_2[179] + mult_out_3[179]) % 3329;
                                                                                                                                                                  mul_add_t[0][180] <= (mult_out_1[180] + mult_out_2[180] + mult_out_3[180]) % 3329;
                                                                                                                                                                  mul_add_t[0][181] <= (mult_out_1[181] + mult_out_2[181] + mult_out_3[181]) % 3329;
                                                                                                                                                                  mul_add_t[0][182] <= (mult_out_1[182] + mult_out_2[182] + mult_out_3[182]) % 3329;
                                                                                                                                                                  mul_add_t[0][183] <= (mult_out_1[183] + mult_out_2[183] + mult_out_3[183]) % 3329;
                                                                                                                                                                  mul_add_t[0][184] <= (mult_out_1[184] + mult_out_2[184] + mult_out_3[184]) % 3329;
                                                                                                                                                                  mul_add_t[0][185] <= (mult_out_1[185] + mult_out_2[185] + mult_out_3[185]) % 3329;
                                                                                                                                                                  mul_add_t[0][186] <= (mult_out_1[186] + mult_out_2[186] + mult_out_3[186]) % 3329;
                                                                                                                                                                  mul_add_t[0][187] <= (mult_out_1[187] + mult_out_2[187] + mult_out_3[187]) % 3329;
                                                                                                                                                                  mul_add_t[0][188] <= (mult_out_1[188] + mult_out_2[188] + mult_out_3[188]) % 3329;
                                                                                                                                                                  mul_add_t[0][189] <= (mult_out_1[189] + mult_out_2[189] + mult_out_3[189]) % 3329;
                                                                                                                                                                  mul_add_t[0][190] <= (mult_out_1[190] + mult_out_2[190] + mult_out_3[190]) % 3329;
                                                                                                                                                                  mul_add_t[0][191] <= (mult_out_1[191] + mult_out_2[191] + mult_out_3[191]) % 3329;
                                                                                                                                                                  mul_add_t[0][192] <= (mult_out_1[192] + mult_out_2[192] + mult_out_3[192]) % 3329;
                                                                                                                                                                  mul_add_t[0][193] <= (mult_out_1[193] + mult_out_2[193] + mult_out_3[193]) % 3329;
                                                                                                                                                                  mul_add_t[0][194] <= (mult_out_1[194] + mult_out_2[194] + mult_out_3[194]) % 3329;
                                                                                                                                                                  mul_add_t[0][195] <= (mult_out_1[195] + mult_out_2[195] + mult_out_3[195]) % 3329;
                                                                                                                                                                  mul_add_t[0][196] <= (mult_out_1[196] + mult_out_2[196] + mult_out_3[196]) % 3329;
                                                                                                                                                                  mul_add_t[0][197] <= (mult_out_1[197] + mult_out_2[197] + mult_out_3[197]) % 3329;
                                                                                                                                                                  mul_add_t[0][198] <= (mult_out_1[198] + mult_out_2[198] + mult_out_3[198]) % 3329;
                                                                                                                                                                  mul_add_t[0][199] <= (mult_out_1[199] + mult_out_2[199] + mult_out_3[199]) % 3329;
                                                                                                                                                                  mul_add_t[0][200] <= (mult_out_1[200] + mult_out_2[200] + mult_out_3[200]) % 3329;
                                                                                                                                                                  mul_add_t[0][201] <= (mult_out_1[201] + mult_out_2[201] + mult_out_3[201]) % 3329;
                                                                                                                                                                  mul_add_t[0][202] <= (mult_out_1[202] + mult_out_2[202] + mult_out_3[202]) % 3329;
                                                                                                                                                                  mul_add_t[0][203] <= (mult_out_1[203] + mult_out_2[203] + mult_out_3[203]) % 3329;
                                                                                                                                                                  mul_add_t[0][204] <= (mult_out_1[204] + mult_out_2[204] + mult_out_3[204]) % 3329;
                                                                                                                                                                  mul_add_t[0][205] <= (mult_out_1[205] + mult_out_2[205] + mult_out_3[205]) % 3329;
                                                                                                                                                                  mul_add_t[0][206] <= (mult_out_1[206] + mult_out_2[206] + mult_out_3[206]) % 3329;
                                                                                                                                                                  mul_add_t[0][207] <= (mult_out_1[207] + mult_out_2[207] + mult_out_3[207]) % 3329;
                                                                                                                                                                  mul_add_t[0][208] <= (mult_out_1[208] + mult_out_2[208] + mult_out_3[208]) % 3329;
                                                                                                                                                                  mul_add_t[0][209] <= (mult_out_1[209] + mult_out_2[209] + mult_out_3[209]) % 3329;
                                                                                                                                                                  mul_add_t[0][210] <= (mult_out_1[210] + mult_out_2[210] + mult_out_3[210]) % 3329;
                                                                                                                                                                  mul_add_t[0][211] <= (mult_out_1[211] + mult_out_2[211] + mult_out_3[211]) % 3329;
                                                                                                                                                                  mul_add_t[0][212] <= (mult_out_1[212] + mult_out_2[212] + mult_out_3[212]) % 3329;
                                                                                                                                                                  mul_add_t[0][213] <= (mult_out_1[213] + mult_out_2[213] + mult_out_3[213]) % 3329;
                                                                                                                                                                  mul_add_t[0][214] <= (mult_out_1[214] + mult_out_2[214] + mult_out_3[214]) % 3329;
                                                                                                                                                                  mul_add_t[0][215] <= (mult_out_1[215] + mult_out_2[215] + mult_out_3[215]) % 3329;
                                                                                                                                                                  mul_add_t[0][216] <= (mult_out_1[216] + mult_out_2[216] + mult_out_3[216]) % 3329;
                                                                                                                                                                  mul_add_t[0][217] <= (mult_out_1[217] + mult_out_2[217] + mult_out_3[217]) % 3329;
                                                                                                                                                                  mul_add_t[0][218] <= (mult_out_1[218] + mult_out_2[218] + mult_out_3[218]) % 3329;
                                                                                                                                                                  mul_add_t[0][219] <= (mult_out_1[219] + mult_out_2[219] + mult_out_3[219]) % 3329;
                                                                                                                                                                  mul_add_t[0][220] <= (mult_out_1[220] + mult_out_2[220] + mult_out_3[220]) % 3329;
                                                                                                                                                                  mul_add_t[0][221] <= (mult_out_1[221] + mult_out_2[221] + mult_out_3[221]) % 3329;
                                                                                                                                                                  mul_add_t[0][222] <= (mult_out_1[222] + mult_out_2[222] + mult_out_3[222]) % 3329;
                                                                                                                                                                  mul_add_t[0][223] <= (mult_out_1[223] + mult_out_2[223] + mult_out_3[223]) % 3329;
                                                                                                                                                                  mul_add_t[0][224] <= (mult_out_1[224] + mult_out_2[224] + mult_out_3[224]) % 3329;
                                                                                                                                                                  mul_add_t[0][225] <= (mult_out_1[225] + mult_out_2[225] + mult_out_3[225]) % 3329;
                                                                                                                                                                  mul_add_t[0][226] <= (mult_out_1[226] + mult_out_2[226] + mult_out_3[226]) % 3329;
                                                                                                                                                                  mul_add_t[0][227] <= (mult_out_1[227] + mult_out_2[227] + mult_out_3[227]) % 3329;
                                                                                                                                                                  mul_add_t[0][228] <= (mult_out_1[228] + mult_out_2[228] + mult_out_3[228]) % 3329;
                                                                                                                                                                  mul_add_t[0][229] <= (mult_out_1[229] + mult_out_2[229] + mult_out_3[229]) % 3329;
                                                                                                                                                                  mul_add_t[0][230] <= (mult_out_1[230] + mult_out_2[230] + mult_out_3[230]) % 3329;
                                                                                                                                                                  mul_add_t[0][231] <= (mult_out_1[231] + mult_out_2[231] + mult_out_3[231]) % 3329;
                                                                                                                                                                  mul_add_t[0][232] <= (mult_out_1[232] + mult_out_2[232] + mult_out_3[232]) % 3329;
                                                                                                                                                                  mul_add_t[0][233] <= (mult_out_1[233] + mult_out_2[233] + mult_out_3[233]) % 3329;
                                                                                                                                                                  mul_add_t[0][234] <= (mult_out_1[234] + mult_out_2[234] + mult_out_3[234]) % 3329;
                                                                                                                                                                  mul_add_t[0][235] <= (mult_out_1[235] + mult_out_2[235] + mult_out_3[235]) % 3329;
                                                                                                                                                                  mul_add_t[0][236] <= (mult_out_1[236] + mult_out_2[236] + mult_out_3[236]) % 3329;
                                                                                                                                                                  mul_add_t[0][237] <= (mult_out_1[237] + mult_out_2[237] + mult_out_3[237]) % 3329;
                                                                                                                                                                  mul_add_t[0][238] <= (mult_out_1[238] + mult_out_2[238] + mult_out_3[238]) % 3329;
                                                                                                                                                                  mul_add_t[0][239] <= (mult_out_1[239] + mult_out_2[239] + mult_out_3[239]) % 3329;
                                                                                                                                                                  mul_add_t[0][240] <= (mult_out_1[240] + mult_out_2[240] + mult_out_3[240]) % 3329;
                                                                                                                                                                  mul_add_t[0][241] <= (mult_out_1[241] + mult_out_2[241] + mult_out_3[241]) % 3329;
                                                                                                                                                                  mul_add_t[0][242] <= (mult_out_1[242] + mult_out_2[242] + mult_out_3[242]) % 3329;
                                                                                                                                                                  mul_add_t[0][243] <= (mult_out_1[243] + mult_out_2[243] + mult_out_3[243]) % 3329;
                                                                                                                                                                  mul_add_t[0][244] <= (mult_out_1[244] + mult_out_2[244] + mult_out_3[244]) % 3329;
                                                                                                                                                                  mul_add_t[0][245] <= (mult_out_1[245] + mult_out_2[245] + mult_out_3[245]) % 3329;
                                                                                                                                                                  mul_add_t[0][246] <= (mult_out_1[246] + mult_out_2[246] + mult_out_3[246]) % 3329;
                                                                                                                                                                  mul_add_t[0][247] <= (mult_out_1[247] + mult_out_2[247] + mult_out_3[247]) % 3329;
                                                                                                                                                                  mul_add_t[0][248] <= (mult_out_1[248] + mult_out_2[248] + mult_out_3[248]) % 3329;
                                                                                                                                                                  mul_add_t[0][249] <= (mult_out_1[249] + mult_out_2[249] + mult_out_3[249]) % 3329;
                                                                                                                                                                  mul_add_t[0][250] <= (mult_out_1[250] + mult_out_2[250] + mult_out_3[250]) % 3329;
                                                                                                                                                                  mul_add_t[0][251] <= (mult_out_1[251] + mult_out_2[251] + mult_out_3[251]) % 3329;
                                                                                                                                                                  mul_add_t[0][252] <= (mult_out_1[252] + mult_out_2[252] + mult_out_3[252]) % 3329;
                                                                                                                                                                  mul_add_t[0][253] <= (mult_out_1[253] + mult_out_2[253] + mult_out_3[253]) % 3329;
                                                                                                                                                                  mul_add_t[0][254] <= (mult_out_1[254] + mult_out_2[254] + mult_out_3[254]) % 3329;
                                                                                                                                                                  mul_add_t[0][255] <= (mult_out_1[255] + mult_out_2[255] + mult_out_3[255]) % 3329;
                                                                                                                                                                   mul_add_t[1][0] <= (mult_out_1[0] + mult_out_2[0] + mult_out_3[0]) % 3329;
                                                                                                                                                                         mul_add_t[1][1] <= (mult_out_1[1] + mult_out_2[1] + mult_out_3[1]) % 3329;
                                                                                                                                                                         mul_add_t[1][2] <= (mult_out_1[2] + mult_out_2[2] + mult_out_3[2]) % 3329;
                                                                                                                                                                         mul_add_t[1][3] <= (mult_out_1[3] + mult_out_2[3] + mult_out_3[3]) % 3329;
                                                                                                                                                                         mul_add_t[1][4] <= (mult_out_1[4] + mult_out_2[4] + mult_out_3[4]) % 3329;
                                                                                                                                                                         mul_add_t[1][5] <= (mult_out_1[5] + mult_out_2[5] + mult_out_3[5]) % 3329;
                                                                                                                                                                         mul_add_t[1][6] <= (mult_out_1[6] + mult_out_2[6] + mult_out_3[6]) % 3329;
                                                                                                                                                                         mul_add_t[1][7] <= (mult_out_1[7] + mult_out_2[7] + mult_out_3[7]) % 3329;
                                                                                                                                                                         mul_add_t[1][8] <= (mult_out_1[8] + mult_out_2[8] + mult_out_3[8]) % 3329;
                                                                                                                                                                         mul_add_t[1][9] <= (mult_out_1[9] + mult_out_2[9] + mult_out_3[9]) % 3329;
                                                                                                                                                                         mul_add_t[1][10] <= (mult_out_1[10] + mult_out_2[10] + mult_out_3[10]) % 3329;
                                                                                                                                                                         mul_add_t[1][11] <= (mult_out_1[11] + mult_out_2[11] + mult_out_3[11]) % 3329;
                                                                                                                                                                         mul_add_t[1][12] <= (mult_out_1[12] + mult_out_2[12] + mult_out_3[12]) % 3329;
                                                                                                                                                                         mul_add_t[1][13] <= (mult_out_1[13] + mult_out_2[13] + mult_out_3[13]) % 3329;
                                                                                                                                                                         mul_add_t[1][14] <= (mult_out_1[14] + mult_out_2[14] + mult_out_3[14]) % 3329;
                                                                                                                                                                         mul_add_t[1][15] <= (mult_out_1[15] + mult_out_2[15] + mult_out_3[15]) % 3329;
                                                                                                                                                                         mul_add_t[1][16] <= (mult_out_1[16] + mult_out_2[16] + mult_out_3[16]) % 3329;
                                                                                                                                                                         mul_add_t[1][17] <= (mult_out_1[17] + mult_out_2[17] + mult_out_3[17]) % 3329;
                                                                                                                                                                         mul_add_t[1][18] <= (mult_out_1[18] + mult_out_2[18] + mult_out_3[18]) % 3329;
                                                                                                                                                                         mul_add_t[1][19] <= (mult_out_1[19] + mult_out_2[19] + mult_out_3[19]) % 3329;
                                                                                                                                                                         mul_add_t[1][20] <= (mult_out_1[20] + mult_out_2[20] + mult_out_3[20]) % 3329;
                                                                                                                                                                         mul_add_t[1][21] <= (mult_out_1[21] + mult_out_2[21] + mult_out_3[21]) % 3329;
                                                                                                                                                                         mul_add_t[1][22] <= (mult_out_1[22] + mult_out_2[22] + mult_out_3[22]) % 3329;
                                                                                                                                                                         mul_add_t[1][23] <= (mult_out_1[23] + mult_out_2[23] + mult_out_3[23]) % 3329;
                                                                                                                                                                         mul_add_t[1][24] <= (mult_out_1[24] + mult_out_2[24] + mult_out_3[24]) % 3329;
                                                                                                                                                                         mul_add_t[1][25] <= (mult_out_1[25] + mult_out_2[25] + mult_out_3[25]) % 3329;
                                                                                                                                                                         mul_add_t[1][26] <= (mult_out_1[26] + mult_out_2[26] + mult_out_3[26]) % 3329;
                                                                                                                                                                         mul_add_t[1][27] <= (mult_out_1[27] + mult_out_2[27] + mult_out_3[27]) % 3329;
                                                                                                                                                                         mul_add_t[1][28] <= (mult_out_1[28] + mult_out_2[28] + mult_out_3[28]) % 3329;
                                                                                                                                                                         mul_add_t[1][29] <= (mult_out_1[29] + mult_out_2[29] + mult_out_3[29]) % 3329;
                                                                                                                                                                         mul_add_t[1][30] <= (mult_out_1[30] + mult_out_2[30] + mult_out_3[30]) % 3329;
                                                                                                                                                                         mul_add_t[1][31] <= (mult_out_1[31] + mult_out_2[31] + mult_out_3[31]) % 3329;
                                                                                                                                                                         mul_add_t[1][32] <= (mult_out_1[32] + mult_out_2[32] + mult_out_3[32]) % 3329;
                                                                                                                                                                         mul_add_t[1][33] <= (mult_out_1[33] + mult_out_2[33] + mult_out_3[33]) % 3329;
                                                                                                                                                                         mul_add_t[1][34] <= (mult_out_1[34] + mult_out_2[34] + mult_out_3[34]) % 3329;
                                                                                                                                                                         mul_add_t[1][35] <= (mult_out_1[35] + mult_out_2[35] + mult_out_3[35]) % 3329;
                                                                                                                                                                         mul_add_t[1][36] <= (mult_out_1[36] + mult_out_2[36] + mult_out_3[36]) % 3329;
                                                                                                                                                                         mul_add_t[1][37] <= (mult_out_1[37] + mult_out_2[37] + mult_out_3[37]) % 3329;
                                                                                                                                                                         mul_add_t[1][38] <= (mult_out_1[38] + mult_out_2[38] + mult_out_3[38]) % 3329;
                                                                                                                                                                         mul_add_t[1][39] <= (mult_out_1[39] + mult_out_2[39] + mult_out_3[39]) % 3329;
                                                                                                                                                                         mul_add_t[1][40] <= (mult_out_1[40] + mult_out_2[40] + mult_out_3[40]) % 3329;
                                                                                                                                                                         mul_add_t[1][41] <= (mult_out_1[41] + mult_out_2[41] + mult_out_3[41]) % 3329;
                                                                                                                                                                         mul_add_t[1][42] <= (mult_out_1[42] + mult_out_2[42] + mult_out_3[42]) % 3329;
                                                                                                                                                                         mul_add_t[1][43] <= (mult_out_1[43] + mult_out_2[43] + mult_out_3[43]) % 3329;
                                                                                                                                                                         mul_add_t[1][44] <= (mult_out_1[44] + mult_out_2[44] + mult_out_3[44]) % 3329;
                                                                                                                                                                         mul_add_t[1][45] <= (mult_out_1[45] + mult_out_2[45] + mult_out_3[45]) % 3329;
                                                                                                                                                                         mul_add_t[1][46] <= (mult_out_1[46] + mult_out_2[46] + mult_out_3[46]) % 3329;
                                                                                                                                                                         mul_add_t[1][47] <= (mult_out_1[47] + mult_out_2[47] + mult_out_3[47]) % 3329;
                                                                                                                                                                         mul_add_t[1][48] <= (mult_out_1[48] + mult_out_2[48] + mult_out_3[48]) % 3329;
                                                                                                                                                                         mul_add_t[1][49] <= (mult_out_1[49] + mult_out_2[49] + mult_out_3[49]) % 3329;
                                                                                                                                                                         mul_add_t[1][50] <= (mult_out_1[50] + mult_out_2[50] + mult_out_3[50]) % 3329;
                                                                                                                                                                         mul_add_t[1][51] <= (mult_out_1[51] + mult_out_2[51] + mult_out_3[51]) % 3329;
                                                                                                                                                                         mul_add_t[1][52] <= (mult_out_1[52] + mult_out_2[52] + mult_out_3[52]) % 3329;
                                                                                                                                                                         mul_add_t[1][53] <= (mult_out_1[53] + mult_out_2[53] + mult_out_3[53]) % 3329;
                                                                                                                                                                         mul_add_t[1][54] <= (mult_out_1[54] + mult_out_2[54] + mult_out_3[54]) % 3329;
                                                                                                                                                                         mul_add_t[1][55] <= (mult_out_1[55] + mult_out_2[55] + mult_out_3[55]) % 3329;
                                                                                                                                                                         mul_add_t[1][56] <= (mult_out_1[56] + mult_out_2[56] + mult_out_3[56]) % 3329;
                                                                                                                                                                         mul_add_t[1][57] <= (mult_out_1[57] + mult_out_2[57] + mult_out_3[57]) % 3329;
                                                                                                                                                                         mul_add_t[1][58] <= (mult_out_1[58] + mult_out_2[58] + mult_out_3[58]) % 3329;
                                                                                                                                                                         mul_add_t[1][59] <= (mult_out_1[59] + mult_out_2[59] + mult_out_3[59]) % 3329;
                                                                                                                                                                         mul_add_t[1][60] <= (mult_out_1[60] + mult_out_2[60] + mult_out_3[60]) % 3329;
                                                                                                                                                                         mul_add_t[1][61] <= (mult_out_1[61] + mult_out_2[61] + mult_out_3[61]) % 3329;
                                                                                                                                                                         mul_add_t[1][62] <= (mult_out_1[62] + mult_out_2[62] + mult_out_3[62]) % 3329;
                                                                                                                                                                         mul_add_t[1][63] <= (mult_out_1[63] + mult_out_2[63] + mult_out_3[63]) % 3329;
                                                                                                                                                                         mul_add_t[1][64] <= (mult_out_1[64] + mult_out_2[64] + mult_out_3[64]) % 3329;
                                                                                                                                                                         mul_add_t[1][65] <= (mult_out_1[65] + mult_out_2[65] + mult_out_3[65]) % 3329;
                                                                                                                                                                         mul_add_t[1][66] <= (mult_out_1[66] + mult_out_2[66] + mult_out_3[66]) % 3329;
                                                                                                                                                                         mul_add_t[1][67] <= (mult_out_1[67] + mult_out_2[67] + mult_out_3[67]) % 3329;
                                                                                                                                                                         mul_add_t[1][68] <= (mult_out_1[68] + mult_out_2[68] + mult_out_3[68]) % 3329;
                                                                                                                                                                         mul_add_t[1][69] <= (mult_out_1[69] + mult_out_2[69] + mult_out_3[69]) % 3329;
                                                                                                                                                                         mul_add_t[1][70] <= (mult_out_1[70] + mult_out_2[70] + mult_out_3[70]) % 3329;
                                                                                                                                                                         mul_add_t[1][71] <= (mult_out_1[71] + mult_out_2[71] + mult_out_3[71]) % 3329;
                                                                                                                                                                         mul_add_t[1][72] <= (mult_out_1[72] + mult_out_2[72] + mult_out_3[72]) % 3329;
                                                                                                                                                                         mul_add_t[1][73] <= (mult_out_1[73] + mult_out_2[73] + mult_out_3[73]) % 3329;
                                                                                                                                                                         mul_add_t[1][74] <= (mult_out_1[74] + mult_out_2[74] + mult_out_3[74]) % 3329;
                                                                                                                                                                         mul_add_t[1][75] <= (mult_out_1[75] + mult_out_2[75] + mult_out_3[75]) % 3329;
                                                                                                                                                                         mul_add_t[1][76] <= (mult_out_1[76] + mult_out_2[76] + mult_out_3[76]) % 3329;
                                                                                                                                                                         mul_add_t[1][77] <= (mult_out_1[77] + mult_out_2[77] + mult_out_3[77]) % 3329;
                                                                                                                                                                         mul_add_t[1][78] <= (mult_out_1[78] + mult_out_2[78] + mult_out_3[78]) % 3329;
                                                                                                                                                                         mul_add_t[1][79] <= (mult_out_1[79] + mult_out_2[79] + mult_out_3[79]) % 3329;
                                                                                                                                                                         mul_add_t[1][80] <= (mult_out_1[80] + mult_out_2[80] + mult_out_3[80]) % 3329;
                                                                                                                                                                         mul_add_t[1][81] <= (mult_out_1[81] + mult_out_2[81] + mult_out_3[81]) % 3329;
                                                                                                                                                                         mul_add_t[1][82] <= (mult_out_1[82] + mult_out_2[82] + mult_out_3[82]) % 3329;
                                                                                                                                                                         mul_add_t[1][83] <= (mult_out_1[83] + mult_out_2[83] + mult_out_3[83]) % 3329;
                                                                                                                                                                         mul_add_t[1][84] <= (mult_out_1[84] + mult_out_2[84] + mult_out_3[84]) % 3329;
                                                                                                                                                                         mul_add_t[1][85] <= (mult_out_1[85] + mult_out_2[85] + mult_out_3[85]) % 3329;
                                                                                                                                                                         mul_add_t[1][86] <= (mult_out_1[86] + mult_out_2[86] + mult_out_3[86]) % 3329;
                                                                                                                                                                         mul_add_t[1][87] <= (mult_out_1[87] + mult_out_2[87] + mult_out_3[87]) % 3329;
                                                                                                                                                                         mul_add_t[1][88] <= (mult_out_1[88] + mult_out_2[88] + mult_out_3[88]) % 3329;
                                                                                                                                                                         mul_add_t[1][89] <= (mult_out_1[89] + mult_out_2[89] + mult_out_3[89]) % 3329;
                                                                                                                                                                         mul_add_t[1][90] <= (mult_out_1[90] + mult_out_2[90] + mult_out_3[90]) % 3329;
                                                                                                                                                                         mul_add_t[1][91] <= (mult_out_1[91] + mult_out_2[91] + mult_out_3[91]) % 3329;
                                                                                                                                                                         mul_add_t[1][92] <= (mult_out_1[92] + mult_out_2[92] + mult_out_3[92]) % 3329;
                                                                                                                                                                         mul_add_t[1][93] <= (mult_out_1[93] + mult_out_2[93] + mult_out_3[93]) % 3329;
                                                                                                                                                                         mul_add_t[1][94] <= (mult_out_1[94] + mult_out_2[94] + mult_out_3[94]) % 3329;
                                                                                                                                                                         mul_add_t[1][95] <= (mult_out_1[95] + mult_out_2[95] + mult_out_3[95]) % 3329;
                                                                                                                                                                         mul_add_t[1][96] <= (mult_out_1[96] + mult_out_2[96] + mult_out_3[96]) % 3329;
                                                                                                                                                                         mul_add_t[1][97] <= (mult_out_1[97] + mult_out_2[97] + mult_out_3[97]) % 3329;
                                                                                                                                                                         mul_add_t[1][98] <= (mult_out_1[98] + mult_out_2[98] + mult_out_3[98]) % 3329;
                                                                                                                                                                         mul_add_t[1][99] <= (mult_out_1[99] + mult_out_2[99] + mult_out_3[99]) % 3329;
                                                                                                                                                                         mul_add_t[1][100] <= (mult_out_1[100] + mult_out_2[100] + mult_out_3[100]) % 3329;
                                                                                                                                                                         mul_add_t[1][101] <= (mult_out_1[101] + mult_out_2[101] + mult_out_3[101]) % 3329;
                                                                                                                                                                         mul_add_t[1][102] <= (mult_out_1[102] + mult_out_2[102] + mult_out_3[102]) % 3329;
                                                                                                                                                                         mul_add_t[1][103] <= (mult_out_1[103] + mult_out_2[103] + mult_out_3[103]) % 3329;
                                                                                                                                                                         mul_add_t[1][104] <= (mult_out_1[104] + mult_out_2[104] + mult_out_3[104]) % 3329;
                                                                                                                                                                         mul_add_t[1][105] <= (mult_out_1[105] + mult_out_2[105] + mult_out_3[105]) % 3329;
                                                                                                                                                                         mul_add_t[1][106] <= (mult_out_1[106] + mult_out_2[106] + mult_out_3[106]) % 3329;
                                                                                                                                                                         mul_add_t[1][107] <= (mult_out_1[107] + mult_out_2[107] + mult_out_3[107]) % 3329;
                                                                                                                                                                         mul_add_t[1][108] <= (mult_out_1[108] + mult_out_2[108] + mult_out_3[108]) % 3329;
                                                                                                                                                                         mul_add_t[1][109] <= (mult_out_1[109] + mult_out_2[109] + mult_out_3[109]) % 3329;
                                                                                                                                                                         mul_add_t[1][110] <= (mult_out_1[110] + mult_out_2[110] + mult_out_3[110]) % 3329;
                                                                                                                                                                         mul_add_t[1][111] <= (mult_out_1[111] + mult_out_2[111] + mult_out_3[111]) % 3329;
                                                                                                                                                                         mul_add_t[1][112] <= (mult_out_1[112] + mult_out_2[112] + mult_out_3[112]) % 3329;
                                                                                                                                                                         mul_add_t[1][113] <= (mult_out_1[113] + mult_out_2[113] + mult_out_3[113]) % 3329;
                                                                                                                                                                         mul_add_t[1][114] <= (mult_out_1[114] + mult_out_2[114] + mult_out_3[114]) % 3329;
                                                                                                                                                                         mul_add_t[1][115] <= (mult_out_1[115] + mult_out_2[115] + mult_out_3[115]) % 3329;
                                                                                                                                                                         mul_add_t[1][116] <= (mult_out_1[116] + mult_out_2[116] + mult_out_3[116]) % 3329;
                                                                                                                                                                         mul_add_t[1][117] <= (mult_out_1[117] + mult_out_2[117] + mult_out_3[117]) % 3329;
                                                                                                                                                                         mul_add_t[1][118] <= (mult_out_1[118] + mult_out_2[118] + mult_out_3[118]) % 3329;
                                                                                                                                                                         mul_add_t[1][119] <= (mult_out_1[119] + mult_out_2[119] + mult_out_3[119]) % 3329;
                                                                                                                                                                         mul_add_t[1][120] <= (mult_out_1[120] + mult_out_2[120] + mult_out_3[120]) % 3329;
                                                                                                                                                                         mul_add_t[1][121] <= (mult_out_1[121] + mult_out_2[121] + mult_out_3[121]) % 3329;
                                                                                                                                                                         mul_add_t[1][122] <= (mult_out_1[122] + mult_out_2[122] + mult_out_3[122]) % 3329;
                                                                                                                                                                         mul_add_t[1][123] <= (mult_out_1[123] + mult_out_2[123] + mult_out_3[123]) % 3329;
                                                                                                                                                                         mul_add_t[1][124] <= (mult_out_1[124] + mult_out_2[124] + mult_out_3[124]) % 3329;
                                                                                                                                                                         mul_add_t[1][125] <= (mult_out_1[125] + mult_out_2[125] + mult_out_3[125]) % 3329;
                                                                                                                                                                         mul_add_t[1][126] <= (mult_out_1[126] + mult_out_2[126] + mult_out_3[126]) % 3329;
                                                                                                                                                                         mul_add_t[1][127] <= (mult_out_1[127] + mult_out_2[127] + mult_out_3[127]) % 3329;
                                                                                                                                                                         mul_add_t[1][128] <= (mult_out_1[128] + mult_out_2[128] + mult_out_3[128]) % 3329;
                                                                                                                                                                         mul_add_t[1][129] <= (mult_out_1[129] + mult_out_2[129] + mult_out_3[129]) % 3329;
                                                                                                                                                                         mul_add_t[1][130] <= (mult_out_1[130] + mult_out_2[130] + mult_out_3[130]) % 3329;
                                                                                                                                                                         mul_add_t[1][131] <= (mult_out_1[131] + mult_out_2[131] + mult_out_3[131]) % 3329;
                                                                                                                                                                         mul_add_t[1][132] <= (mult_out_1[132] + mult_out_2[132] + mult_out_3[132]) % 3329;
                                                                                                                                                                         mul_add_t[1][133] <= (mult_out_1[133] + mult_out_2[133] + mult_out_3[133]) % 3329;
                                                                                                                                                                         mul_add_t[1][134] <= (mult_out_1[134] + mult_out_2[134] + mult_out_3[134]) % 3329;
                                                                                                                                                                         mul_add_t[1][135] <= (mult_out_1[135] + mult_out_2[135] + mult_out_3[135]) % 3329;
                                                                                                                                                                         mul_add_t[1][136] <= (mult_out_1[136] + mult_out_2[136] + mult_out_3[136]) % 3329;
                                                                                                                                                                         mul_add_t[1][137] <= (mult_out_1[137] + mult_out_2[137] + mult_out_3[137]) % 3329;
                                                                                                                                                                         mul_add_t[1][138] <= (mult_out_1[138] + mult_out_2[138] + mult_out_3[138]) % 3329;
                                                                                                                                                                         mul_add_t[1][139] <= (mult_out_1[139] + mult_out_2[139] + mult_out_3[139]) % 3329;
                                                                                                                                                                         mul_add_t[1][140] <= (mult_out_1[140] + mult_out_2[140] + mult_out_3[140]) % 3329;
                                                                                                                                                                         mul_add_t[1][141] <= (mult_out_1[141] + mult_out_2[141] + mult_out_3[141]) % 3329;
                                                                                                                                                                         mul_add_t[1][142] <= (mult_out_1[142] + mult_out_2[142] + mult_out_3[142]) % 3329;
                                                                                                                                                                         mul_add_t[1][143] <= (mult_out_1[143] + mult_out_2[143] + mult_out_3[143]) % 3329;
                                                                                                                                                                         mul_add_t[1][144] <= (mult_out_1[144] + mult_out_2[144] + mult_out_3[144]) % 3329;
                                                                                                                                                                         mul_add_t[1][145] <= (mult_out_1[145] + mult_out_2[145] + mult_out_3[145]) % 3329;
                                                                                                                                                                         mul_add_t[1][146] <= (mult_out_1[146] + mult_out_2[146] + mult_out_3[146]) % 3329;
                                                                                                                                                                         mul_add_t[1][147] <= (mult_out_1[147] + mult_out_2[147] + mult_out_3[147]) % 3329;
                                                                                                                                                                         mul_add_t[1][148] <= (mult_out_1[148] + mult_out_2[148] + mult_out_3[148]) % 3329;
                                                                                                                                                                         mul_add_t[1][149] <= (mult_out_1[149] + mult_out_2[149] + mult_out_3[149]) % 3329;
                                                                                                                                                                         mul_add_t[1][150] <= (mult_out_1[150] + mult_out_2[150] + mult_out_3[150]) % 3329;
                                                                                                                                                                         mul_add_t[1][151] <= (mult_out_1[151] + mult_out_2[151] + mult_out_3[151]) % 3329;
                                                                                                                                                                         mul_add_t[1][152] <= (mult_out_1[152] + mult_out_2[152] + mult_out_3[152]) % 3329;
                                                                                                                                                                         mul_add_t[1][153] <= (mult_out_1[153] + mult_out_2[153] + mult_out_3[153]) % 3329;
                                                                                                                                                                         mul_add_t[1][154] <= (mult_out_1[154] + mult_out_2[154] + mult_out_3[154]) % 3329;
                                                                                                                                                                         mul_add_t[1][155] <= (mult_out_1[155] + mult_out_2[155] + mult_out_3[155]) % 3329;
                                                                                                                                                                         mul_add_t[1][156] <= (mult_out_1[156] + mult_out_2[156] + mult_out_3[156]) % 3329;
                                                                                                                                                                         mul_add_t[1][157] <= (mult_out_1[157] + mult_out_2[157] + mult_out_3[157]) % 3329;
                                                                                                                                                                         mul_add_t[1][158] <= (mult_out_1[158] + mult_out_2[158] + mult_out_3[158]) % 3329;
                                                                                                                                                                         mul_add_t[1][159] <= (mult_out_1[159] + mult_out_2[159] + mult_out_3[159]) % 3329;
                                                                                                                                                                         mul_add_t[1][160] <= (mult_out_1[160] + mult_out_2[160] + mult_out_3[160]) % 3329;
                                                                                                                                                                         mul_add_t[1][161] <= (mult_out_1[161] + mult_out_2[161] + mult_out_3[161]) % 3329;
                                                                                                                                                                         mul_add_t[1][162] <= (mult_out_1[162] + mult_out_2[162] + mult_out_3[162]) % 3329;
                                                                                                                                                                         mul_add_t[1][163] <= (mult_out_1[163] + mult_out_2[163] + mult_out_3[163]) % 3329;
                                                                                                                                                                         mul_add_t[1][164] <= (mult_out_1[164] + mult_out_2[164] + mult_out_3[164]) % 3329;
                                                                                                                                                                         mul_add_t[1][165] <= (mult_out_1[165] + mult_out_2[165] + mult_out_3[165]) % 3329;
                                                                                                                                                                         mul_add_t[1][166] <= (mult_out_1[166] + mult_out_2[166] + mult_out_3[166]) % 3329;
                                                                                                                                                                         mul_add_t[1][167] <= (mult_out_1[167] + mult_out_2[167] + mult_out_3[167]) % 3329;
                                                                                                                                                                         mul_add_t[1][168] <= (mult_out_1[168] + mult_out_2[168] + mult_out_3[168]) % 3329;
                                                                                                                                                                         mul_add_t[1][169] <= (mult_out_1[169] + mult_out_2[169] + mult_out_3[169]) % 3329;
                                                                                                                                                                         mul_add_t[1][170] <= (mult_out_1[170] + mult_out_2[170] + mult_out_3[170]) % 3329;
                                                                                                                                                                         mul_add_t[1][171] <= (mult_out_1[171] + mult_out_2[171] + mult_out_3[171]) % 3329;
                                                                                                                                                                         mul_add_t[1][172] <= (mult_out_1[172] + mult_out_2[172] + mult_out_3[172]) % 3329;
                                                                                                                                                                         mul_add_t[1][173] <= (mult_out_1[173] + mult_out_2[173] + mult_out_3[173]) % 3329;
                                                                                                                                                                         mul_add_t[1][174] <= (mult_out_1[174] + mult_out_2[174] + mult_out_3[174]) % 3329;
                                                                                                                                                                         mul_add_t[1][175] <= (mult_out_1[175] + mult_out_2[175] + mult_out_3[175]) % 3329;
                                                                                                                                                                         mul_add_t[1][176] <= (mult_out_1[176] + mult_out_2[176] + mult_out_3[176]) % 3329;
                                                                                                                                                                         mul_add_t[1][177] <= (mult_out_1[177] + mult_out_2[177] + mult_out_3[177]) % 3329;
                                                                                                                                                                         mul_add_t[1][178] <= (mult_out_1[178] + mult_out_2[178] + mult_out_3[178]) % 3329;
                                                                                                                                                                         mul_add_t[1][179] <= (mult_out_1[179] + mult_out_2[179] + mult_out_3[179]) % 3329;
                                                                                                                                                                         mul_add_t[1][180] <= (mult_out_1[180] + mult_out_2[180] + mult_out_3[180]) % 3329;
                                                                                                                                                                         mul_add_t[1][181] <= (mult_out_1[181] + mult_out_2[181] + mult_out_3[181]) % 3329;
                                                                                                                                                                         mul_add_t[1][182] <= (mult_out_1[182] + mult_out_2[182] + mult_out_3[182]) % 3329;
                                                                                                                                                                         mul_add_t[1][183] <= (mult_out_1[183] + mult_out_2[183] + mult_out_3[183]) % 3329;
                                                                                                                                                                         mul_add_t[1][184] <= (mult_out_1[184] + mult_out_2[184] + mult_out_3[184]) % 3329;
                                                                                                                                                                         mul_add_t[1][185] <= (mult_out_1[185] + mult_out_2[185] + mult_out_3[185]) % 3329;
                                                                                                                                                                         mul_add_t[1][186] <= (mult_out_1[186] + mult_out_2[186] + mult_out_3[186]) % 3329;
                                                                                                                                                                         mul_add_t[1][187] <= (mult_out_1[187] + mult_out_2[187] + mult_out_3[187]) % 3329;
                                                                                                                                                                         mul_add_t[1][188] <= (mult_out_1[188] + mult_out_2[188] + mult_out_3[188]) % 3329;
                                                                                                                                                                         mul_add_t[1][189] <= (mult_out_1[189] + mult_out_2[189] + mult_out_3[189]) % 3329;
                                                                                                                                                                         mul_add_t[1][190] <= (mult_out_1[190] + mult_out_2[190] + mult_out_3[190]) % 3329;
                                                                                                                                                                         mul_add_t[1][191] <= (mult_out_1[191] + mult_out_2[191] + mult_out_3[191]) % 3329;
                                                                                                                                                                         mul_add_t[1][192] <= (mult_out_1[192] + mult_out_2[192] + mult_out_3[192]) % 3329;
                                                                                                                                                                         mul_add_t[1][193] <= (mult_out_1[193] + mult_out_2[193] + mult_out_3[193]) % 3329;
                                                                                                                                                                         mul_add_t[1][194] <= (mult_out_1[194] + mult_out_2[194] + mult_out_3[194]) % 3329;
                                                                                                                                                                         mul_add_t[1][195] <= (mult_out_1[195] + mult_out_2[195] + mult_out_3[195]) % 3329;
                                                                                                                                                                         mul_add_t[1][196] <= (mult_out_1[196] + mult_out_2[196] + mult_out_3[196]) % 3329;
                                                                                                                                                                         mul_add_t[1][197] <= (mult_out_1[197] + mult_out_2[197] + mult_out_3[197]) % 3329;
                                                                                                                                                                         mul_add_t[1][198] <= (mult_out_1[198] + mult_out_2[198] + mult_out_3[198]) % 3329;
                                                                                                                                                                         mul_add_t[1][199] <= (mult_out_1[199] + mult_out_2[199] + mult_out_3[199]) % 3329;
                                                                                                                                                                         mul_add_t[1][200] <= (mult_out_1[200] + mult_out_2[200] + mult_out_3[200]) % 3329;
                                                                                                                                                                         mul_add_t[1][201] <= (mult_out_1[201] + mult_out_2[201] + mult_out_3[201]) % 3329;
                                                                                                                                                                         mul_add_t[1][202] <= (mult_out_1[202] + mult_out_2[202] + mult_out_3[202]) % 3329;
                                                                                                                                                                         mul_add_t[1][203] <= (mult_out_1[203] + mult_out_2[203] + mult_out_3[203]) % 3329;
                                                                                                                                                                         mul_add_t[1][204] <= (mult_out_1[204] + mult_out_2[204] + mult_out_3[204]) % 3329;
                                                                                                                                                                         mul_add_t[1][205] <= (mult_out_1[205] + mult_out_2[205] + mult_out_3[205]) % 3329;
                                                                                                                                                                         mul_add_t[1][206] <= (mult_out_1[206] + mult_out_2[206] + mult_out_3[206]) % 3329;
                                                                                                                                                                         mul_add_t[1][207] <= (mult_out_1[207] + mult_out_2[207] + mult_out_3[207]) % 3329;
                                                                                                                                                                         mul_add_t[1][208] <= (mult_out_1[208] + mult_out_2[208] + mult_out_3[208]) % 3329;
                                                                                                                                                                         mul_add_t[1][209] <= (mult_out_1[209] + mult_out_2[209] + mult_out_3[209]) % 3329;
                                                                                                                                                                         mul_add_t[1][210] <= (mult_out_1[210] + mult_out_2[210] + mult_out_3[210]) % 3329;
                                                                                                                                                                         mul_add_t[1][211] <= (mult_out_1[211] + mult_out_2[211] + mult_out_3[211]) % 3329;
                                                                                                                                                                         mul_add_t[1][212] <= (mult_out_1[212] + mult_out_2[212] + mult_out_3[212]) % 3329;
                                                                                                                                                                         mul_add_t[1][213] <= (mult_out_1[213] + mult_out_2[213] + mult_out_3[213]) % 3329;
                                                                                                                                                                         mul_add_t[1][214] <= (mult_out_1[214] + mult_out_2[214] + mult_out_3[214]) % 3329;
                                                                                                                                                                         mul_add_t[1][215] <= (mult_out_1[215] + mult_out_2[215] + mult_out_3[215]) % 3329;
                                                                                                                                                                         mul_add_t[1][216] <= (mult_out_1[216] + mult_out_2[216] + mult_out_3[216]) % 3329;
                                                                                                                                                                         mul_add_t[1][217] <= (mult_out_1[217] + mult_out_2[217] + mult_out_3[217]) % 3329;
                                                                                                                                                                         mul_add_t[1][218] <= (mult_out_1[218] + mult_out_2[218] + mult_out_3[218]) % 3329;
                                                                                                                                                                         mul_add_t[1][219] <= (mult_out_1[219] + mult_out_2[219] + mult_out_3[219]) % 3329;
                                                                                                                                                                         mul_add_t[1][220] <= (mult_out_1[220] + mult_out_2[220] + mult_out_3[220]) % 3329;
                                                                                                                                                                         mul_add_t[1][221] <= (mult_out_1[221] + mult_out_2[221] + mult_out_3[221]) % 3329;
                                                                                                                                                                         mul_add_t[1][222] <= (mult_out_1[222] + mult_out_2[222] + mult_out_3[222]) % 3329;
                                                                                                                                                                         mul_add_t[1][223] <= (mult_out_1[223] + mult_out_2[223] + mult_out_3[223]) % 3329;
                                                                                                                                                                         mul_add_t[1][224] <= (mult_out_1[224] + mult_out_2[224] + mult_out_3[224]) % 3329;
                                                                                                                                                                         mul_add_t[1][225] <= (mult_out_1[225] + mult_out_2[225] + mult_out_3[225]) % 3329;
                                                                                                                                                                         mul_add_t[1][226] <= (mult_out_1[226] + mult_out_2[226] + mult_out_3[226]) % 3329;
                                                                                                                                                                         mul_add_t[1][227] <= (mult_out_1[227] + mult_out_2[227] + mult_out_3[227]) % 3329;
                                                                                                                                                                         mul_add_t[1][228] <= (mult_out_1[228] + mult_out_2[228] + mult_out_3[228]) % 3329;
                                                                                                                                                                         mul_add_t[1][229] <= (mult_out_1[229] + mult_out_2[229] + mult_out_3[229]) % 3329;
                                                                                                                                                                         mul_add_t[1][230] <= (mult_out_1[230] + mult_out_2[230] + mult_out_3[230]) % 3329;
                                                                                                                                                                         mul_add_t[1][231] <= (mult_out_1[231] + mult_out_2[231] + mult_out_3[231]) % 3329;
                                                                                                                                                                         mul_add_t[1][232] <= (mult_out_1[232] + mult_out_2[232] + mult_out_3[232]) % 3329;
                                                                                                                                                                         mul_add_t[1][233] <= (mult_out_1[233] + mult_out_2[233] + mult_out_3[233]) % 3329;
                                                                                                                                                                         mul_add_t[1][234] <= (mult_out_1[234] + mult_out_2[234] + mult_out_3[234]) % 3329;
                                                                                                                                                                         mul_add_t[1][235] <= (mult_out_1[235] + mult_out_2[235] + mult_out_3[235]) % 3329;
                                                                                                                                                                         mul_add_t[1][236] <= (mult_out_1[236] + mult_out_2[236] + mult_out_3[236]) % 3329;
                                                                                                                                                                         mul_add_t[1][237] <= (mult_out_1[237] + mult_out_2[237] + mult_out_3[237]) % 3329;
                                                                                                                                                                         mul_add_t[1][238] <= (mult_out_1[238] + mult_out_2[238] + mult_out_3[238]) % 3329;
                                                                                                                                                                         mul_add_t[1][239] <= (mult_out_1[239] + mult_out_2[239] + mult_out_3[239]) % 3329;
                                                                                                                                                                         mul_add_t[1][240] <= (mult_out_1[240] + mult_out_2[240] + mult_out_3[240]) % 3329;
                                                                                                                                                                         mul_add_t[1][241] <= (mult_out_1[241] + mult_out_2[241] + mult_out_3[241]) % 3329;
                                                                                                                                                                         mul_add_t[1][242] <= (mult_out_1[242] + mult_out_2[242] + mult_out_3[242]) % 3329;
                                                                                                                                                                         mul_add_t[1][243] <= (mult_out_1[243] + mult_out_2[243] + mult_out_3[243]) % 3329;
                                                                                                                                                                         mul_add_t[1][244] <= (mult_out_1[244] + mult_out_2[244] + mult_out_3[244]) % 3329;
                                                                                                                                                                         mul_add_t[1][245] <= (mult_out_1[245] + mult_out_2[245] + mult_out_3[245]) % 3329;
                                                                                                                                                                         mul_add_t[1][246] <= (mult_out_1[246] + mult_out_2[246] + mult_out_3[246]) % 3329;
                                                                                                                                                                         mul_add_t[1][247] <= (mult_out_1[247] + mult_out_2[247] + mult_out_3[247]) % 3329;
                                                                                                                                                                         mul_add_t[1][248] <= (mult_out_1[248] + mult_out_2[248] + mult_out_3[248]) % 3329;
                                                                                                                                                                         mul_add_t[1][249] <= (mult_out_1[249] + mult_out_2[249] + mult_out_3[249]) % 3329;
                                                                                                                                                                         mul_add_t[1][250] <= (mult_out_1[250] + mult_out_2[250] + mult_out_3[250]) % 3329;
                                                                                                                                                                         mul_add_t[1][251] <= (mult_out_1[251] + mult_out_2[251] + mult_out_3[251]) % 3329;
                                                                                                                                                                         mul_add_t[1][252] <= (mult_out_1[252] + mult_out_2[252] + mult_out_3[252]) % 3329;
                                                                                                                                                                         mul_add_t[1][253] <= (mult_out_1[253] + mult_out_2[253] + mult_out_3[253]) % 3329;
                                                                                                                                                                         mul_add_t[1][254] <= (mult_out_1[254] + mult_out_2[254] + mult_out_3[254]) % 3329;
                                                                                                                                                                         mul_add_t[1][255] <= (mult_out_1[255] + mult_out_2[255] + mult_out_3[255]) % 3329;
                                                                                                                                                                         mul_add_t[2][0] <= (mult_out_1[0] + mult_out_2[0] + mult_out_3[0]) % 3329;
                                                                                                                                                                                 mul_add_t[2][1] <= (mult_out_1[1] + mult_out_2[1] + mult_out_3[1]) % 3329;
                                                                                                                                                                                 mul_add_t[2][2] <= (mult_out_1[2] + mult_out_2[2] + mult_out_3[2]) % 3329;
                                                                                                                                                                                 mul_add_t[2][3] <= (mult_out_1[3] + mult_out_2[3] + mult_out_3[3]) % 3329;
                                                                                                                                                                                 mul_add_t[2][4] <= (mult_out_1[4] + mult_out_2[4] + mult_out_3[4]) % 3329;
                                                                                                                                                                                 mul_add_t[2][5] <= (mult_out_1[5] + mult_out_2[5] + mult_out_3[5]) % 3329;
                                                                                                                                                                                 mul_add_t[2][6] <= (mult_out_1[6] + mult_out_2[6] + mult_out_3[6]) % 3329;
                                                                                                                                                                                 mul_add_t[2][7] <= (mult_out_1[7] + mult_out_2[7] + mult_out_3[7]) % 3329;
                                                                                                                                                                                 mul_add_t[2][8] <= (mult_out_1[8] + mult_out_2[8] + mult_out_3[8]) % 3329;
                                                                                                                                                                                 mul_add_t[2][9] <= (mult_out_1[9] + mult_out_2[9] + mult_out_3[9]) % 3329;
                                                                                                                                                                                 mul_add_t[2][10] <= (mult_out_1[10] + mult_out_2[10] + mult_out_3[10]) % 3329;
                                                                                                                                                                                 mul_add_t[2][11] <= (mult_out_1[11] + mult_out_2[11] + mult_out_3[11]) % 3329;
                                                                                                                                                                                 mul_add_t[2][12] <= (mult_out_1[12] + mult_out_2[12] + mult_out_3[12]) % 3329;
                                                                                                                                                                                 mul_add_t[2][13] <= (mult_out_1[13] + mult_out_2[13] + mult_out_3[13]) % 3329;
                                                                                                                                                                                 mul_add_t[2][14] <= (mult_out_1[14] + mult_out_2[14] + mult_out_3[14]) % 3329;
                                                                                                                                                                                 mul_add_t[2][15] <= (mult_out_1[15] + mult_out_2[15] + mult_out_3[15]) % 3329;
                                                                                                                                                                                 mul_add_t[2][16] <= (mult_out_1[16] + mult_out_2[16] + mult_out_3[16]) % 3329;
                                                                                                                                                                                 mul_add_t[2][17] <= (mult_out_1[17] + mult_out_2[17] + mult_out_3[17]) % 3329;
                                                                                                                                                                                 mul_add_t[2][18] <= (mult_out_1[18] + mult_out_2[18] + mult_out_3[18]) % 3329;
                                                                                                                                                                                 mul_add_t[2][19] <= (mult_out_1[19] + mult_out_2[19] + mult_out_3[19]) % 3329;
                                                                                                                                                                                 mul_add_t[2][20] <= (mult_out_1[20] + mult_out_2[20] + mult_out_3[20]) % 3329;
                                                                                                                                                                                 mul_add_t[2][21] <= (mult_out_1[21] + mult_out_2[21] + mult_out_3[21]) % 3329;
                                                                                                                                                                                 mul_add_t[2][22] <= (mult_out_1[22] + mult_out_2[22] + mult_out_3[22]) % 3329;
                                                                                                                                                                                 mul_add_t[2][23] <= (mult_out_1[23] + mult_out_2[23] + mult_out_3[23]) % 3329;
                                                                                                                                                                                 mul_add_t[2][24] <= (mult_out_1[24] + mult_out_2[24] + mult_out_3[24]) % 3329;
                                                                                                                                                                                 mul_add_t[2][25] <= (mult_out_1[25] + mult_out_2[25] + mult_out_3[25]) % 3329;
                                                                                                                                                                                 mul_add_t[2][26] <= (mult_out_1[26] + mult_out_2[26] + mult_out_3[26]) % 3329;
                                                                                                                                                                                 mul_add_t[2][27] <= (mult_out_1[27] + mult_out_2[27] + mult_out_3[27]) % 3329;
                                                                                                                                                                                 mul_add_t[2][28] <= (mult_out_1[28] + mult_out_2[28] + mult_out_3[28]) % 3329;
                                                                                                                                                                                 mul_add_t[2][29] <= (mult_out_1[29] + mult_out_2[29] + mult_out_3[29]) % 3329;
                                                                                                                                                                                 mul_add_t[2][30] <= (mult_out_1[30] + mult_out_2[30] + mult_out_3[30]) % 3329;
                                                                                                                                                                                 mul_add_t[2][31] <= (mult_out_1[31] + mult_out_2[31] + mult_out_3[31]) % 3329;
                                                                                                                                                                                 mul_add_t[2][32] <= (mult_out_1[32] + mult_out_2[32] + mult_out_3[32]) % 3329;
                                                                                                                                                                                 mul_add_t[2][33] <= (mult_out_1[33] + mult_out_2[33] + mult_out_3[33]) % 3329;
                                                                                                                                                                                 mul_add_t[2][34] <= (mult_out_1[34] + mult_out_2[34] + mult_out_3[34]) % 3329;
                                                                                                                                                                                 mul_add_t[2][35] <= (mult_out_1[35] + mult_out_2[35] + mult_out_3[35]) % 3329;
                                                                                                                                                                                 mul_add_t[2][36] <= (mult_out_1[36] + mult_out_2[36] + mult_out_3[36]) % 3329;
                                                                                                                                                                                 mul_add_t[2][37] <= (mult_out_1[37] + mult_out_2[37] + mult_out_3[37]) % 3329;
                                                                                                                                                                                 mul_add_t[2][38] <= (mult_out_1[38] + mult_out_2[38] + mult_out_3[38]) % 3329;
                                                                                                                                                                                 mul_add_t[2][39] <= (mult_out_1[39] + mult_out_2[39] + mult_out_3[39]) % 3329;
                                                                                                                                                                                 mul_add_t[2][40] <= (mult_out_1[40] + mult_out_2[40] + mult_out_3[40]) % 3329;
                                                                                                                                                                                 mul_add_t[2][41] <= (mult_out_1[41] + mult_out_2[41] + mult_out_3[41]) % 3329;
                                                                                                                                                                                 mul_add_t[2][42] <= (mult_out_1[42] + mult_out_2[42] + mult_out_3[42]) % 3329;
                                                                                                                                                                                 mul_add_t[2][43] <= (mult_out_1[43] + mult_out_2[43] + mult_out_3[43]) % 3329;
                                                                                                                                                                                 mul_add_t[2][44] <= (mult_out_1[44] + mult_out_2[44] + mult_out_3[44]) % 3329;
                                                                                                                                                                                 mul_add_t[2][45] <= (mult_out_1[45] + mult_out_2[45] + mult_out_3[45]) % 3329;
                                                                                                                                                                                 mul_add_t[2][46] <= (mult_out_1[46] + mult_out_2[46] + mult_out_3[46]) % 3329;
                                                                                                                                                                                 mul_add_t[2][47] <= (mult_out_1[47] + mult_out_2[47] + mult_out_3[47]) % 3329;
                                                                                                                                                                                 mul_add_t[2][48] <= (mult_out_1[48] + mult_out_2[48] + mult_out_3[48]) % 3329;
                                                                                                                                                                                 mul_add_t[2][49] <= (mult_out_1[49] + mult_out_2[49] + mult_out_3[49]) % 3329;
                                                                                                                                                                                 mul_add_t[2][50] <= (mult_out_1[50] + mult_out_2[50] + mult_out_3[50]) % 3329;
                                                                                                                                                                                 mul_add_t[2][51] <= (mult_out_1[51] + mult_out_2[51] + mult_out_3[51]) % 3329;
                                                                                                                                                                                 mul_add_t[2][52] <= (mult_out_1[52] + mult_out_2[52] + mult_out_3[52]) % 3329;
                                                                                                                                                                                 mul_add_t[2][53] <= (mult_out_1[53] + mult_out_2[53] + mult_out_3[53]) % 3329;
                                                                                                                                                                                 mul_add_t[2][54] <= (mult_out_1[54] + mult_out_2[54] + mult_out_3[54]) % 3329;
                                                                                                                                                                                 mul_add_t[2][55] <= (mult_out_1[55] + mult_out_2[55] + mult_out_3[55]) % 3329;
                                                                                                                                                                                 mul_add_t[2][56] <= (mult_out_1[56] + mult_out_2[56] + mult_out_3[56]) % 3329;
                                                                                                                                                                                 mul_add_t[2][57] <= (mult_out_1[57] + mult_out_2[57] + mult_out_3[57]) % 3329;
                                                                                                                                                                                 mul_add_t[2][58] <= (mult_out_1[58] + mult_out_2[58] + mult_out_3[58]) % 3329;
                                                                                                                                                                                 mul_add_t[2][59] <= (mult_out_1[59] + mult_out_2[59] + mult_out_3[59]) % 3329;
                                                                                                                                                                                 mul_add_t[2][60] <= (mult_out_1[60] + mult_out_2[60] + mult_out_3[60]) % 3329;
                                                                                                                                                                                 mul_add_t[2][61] <= (mult_out_1[61] + mult_out_2[61] + mult_out_3[61]) % 3329;
                                                                                                                                                                                 mul_add_t[2][62] <= (mult_out_1[62] + mult_out_2[62] + mult_out_3[62]) % 3329;
                                                                                                                                                                                 mul_add_t[2][63] <= (mult_out_1[63] + mult_out_2[63] + mult_out_3[63]) % 3329;
                                                                                                                                                                                 mul_add_t[2][64] <= (mult_out_1[64] + mult_out_2[64] + mult_out_3[64]) % 3329;
                                                                                                                                                                                 mul_add_t[2][65] <= (mult_out_1[65] + mult_out_2[65] + mult_out_3[65]) % 3329;
                                                                                                                                                                                 mul_add_t[2][66] <= (mult_out_1[66] + mult_out_2[66] + mult_out_3[66]) % 3329;
                                                                                                                                                                                 mul_add_t[2][67] <= (mult_out_1[67] + mult_out_2[67] + mult_out_3[67]) % 3329;
                                                                                                                                                                                 mul_add_t[2][68] <= (mult_out_1[68] + mult_out_2[68] + mult_out_3[68]) % 3329;
                                                                                                                                                                                 mul_add_t[2][69] <= (mult_out_1[69] + mult_out_2[69] + mult_out_3[69]) % 3329;
                                                                                                                                                                                 mul_add_t[2][70] <= (mult_out_1[70] + mult_out_2[70] + mult_out_3[70]) % 3329;
                                                                                                                                                                                 mul_add_t[2][71] <= (mult_out_1[71] + mult_out_2[71] + mult_out_3[71]) % 3329;
                                                                                                                                                                                 mul_add_t[2][72] <= (mult_out_1[72] + mult_out_2[72] + mult_out_3[72]) % 3329;
                                                                                                                                                                                 mul_add_t[2][73] <= (mult_out_1[73] + mult_out_2[73] + mult_out_3[73]) % 3329;
                                                                                                                                                                                 mul_add_t[2][74] <= (mult_out_1[74] + mult_out_2[74] + mult_out_3[74]) % 3329;
                                                                                                                                                                                 mul_add_t[2][75] <= (mult_out_1[75] + mult_out_2[75] + mult_out_3[75]) % 3329;
                                                                                                                                                                                 mul_add_t[2][76] <= (mult_out_1[76] + mult_out_2[76] + mult_out_3[76]) % 3329;
                                                                                                                                                                                 mul_add_t[2][77] <= (mult_out_1[77] + mult_out_2[77] + mult_out_3[77]) % 3329;
                                                                                                                                                                                 mul_add_t[2][78] <= (mult_out_1[78] + mult_out_2[78] + mult_out_3[78]) % 3329;
                                                                                                                                                                                 mul_add_t[2][79] <= (mult_out_1[79] + mult_out_2[79] + mult_out_3[79]) % 3329;
                                                                                                                                                                                 mul_add_t[2][80] <= (mult_out_1[80] + mult_out_2[80] + mult_out_3[80]) % 3329;
                                                                                                                                                                                 mul_add_t[2][81] <= (mult_out_1[81] + mult_out_2[81] + mult_out_3[81]) % 3329;
                                                                                                                                                                                 mul_add_t[2][82] <= (mult_out_1[82] + mult_out_2[82] + mult_out_3[82]) % 3329;
                                                                                                                                                                                 mul_add_t[2][83] <= (mult_out_1[83] + mult_out_2[83] + mult_out_3[83]) % 3329;
                                                                                                                                                                                 mul_add_t[2][84] <= (mult_out_1[84] + mult_out_2[84] + mult_out_3[84]) % 3329;
                                                                                                                                                                                 mul_add_t[2][85] <= (mult_out_1[85] + mult_out_2[85] + mult_out_3[85]) % 3329;
                                                                                                                                                                                 mul_add_t[2][86] <= (mult_out_1[86] + mult_out_2[86] + mult_out_3[86]) % 3329;
                                                                                                                                                                                 mul_add_t[2][87] <= (mult_out_1[87] + mult_out_2[87] + mult_out_3[87]) % 3329;
                                                                                                                                                                                 mul_add_t[2][88] <= (mult_out_1[88] + mult_out_2[88] + mult_out_3[88]) % 3329;
                                                                                                                                                                                 mul_add_t[2][89] <= (mult_out_1[89] + mult_out_2[89] + mult_out_3[89]) % 3329;
                                                                                                                                                                                 mul_add_t[2][90] <= (mult_out_1[90] + mult_out_2[90] + mult_out_3[90]) % 3329;
                                                                                                                                                                                 mul_add_t[2][91] <= (mult_out_1[91] + mult_out_2[91] + mult_out_3[91]) % 3329;
                                                                                                                                                                                 mul_add_t[2][92] <= (mult_out_1[92] + mult_out_2[92] + mult_out_3[92]) % 3329;
                                                                                                                                                                                 mul_add_t[2][93] <= (mult_out_1[93] + mult_out_2[93] + mult_out_3[93]) % 3329;
                                                                                                                                                                                 mul_add_t[2][94] <= (mult_out_1[94] + mult_out_2[94] + mult_out_3[94]) % 3329;
                                                                                                                                                                                 mul_add_t[2][95] <= (mult_out_1[95] + mult_out_2[95] + mult_out_3[95]) % 3329;
                                                                                                                                                                                 mul_add_t[2][96] <= (mult_out_1[96] + mult_out_2[96] + mult_out_3[96]) % 3329;
                                                                                                                                                                                 mul_add_t[2][97] <= (mult_out_1[97] + mult_out_2[97] + mult_out_3[97]) % 3329;
                                                                                                                                                                                 mul_add_t[2][98] <= (mult_out_1[98] + mult_out_2[98] + mult_out_3[98]) % 3329;
                                                                                                                                                                                 mul_add_t[2][99] <= (mult_out_1[99] + mult_out_2[99] + mult_out_3[99]) % 3329;
                                                                                                                                                                                 mul_add_t[2][100] <= (mult_out_1[100] + mult_out_2[100] + mult_out_3[100]) % 3329;
                                                                                                                                                                                 mul_add_t[2][101] <= (mult_out_1[101] + mult_out_2[101] + mult_out_3[101]) % 3329;
                                                                                                                                                                                 mul_add_t[2][102] <= (mult_out_1[102] + mult_out_2[102] + mult_out_3[102]) % 3329;
                                                                                                                                                                                 mul_add_t[2][103] <= (mult_out_1[103] + mult_out_2[103] + mult_out_3[103]) % 3329;
                                                                                                                                                                                 mul_add_t[2][104] <= (mult_out_1[104] + mult_out_2[104] + mult_out_3[104]) % 3329;
                                                                                                                                                                                 mul_add_t[2][105] <= (mult_out_1[105] + mult_out_2[105] + mult_out_3[105]) % 3329;
                                                                                                                                                                                 mul_add_t[2][106] <= (mult_out_1[106] + mult_out_2[106] + mult_out_3[106]) % 3329;
                                                                                                                                                                                 mul_add_t[2][107] <= (mult_out_1[107] + mult_out_2[107] + mult_out_3[107]) % 3329;
                                                                                                                                                                                 mul_add_t[2][108] <= (mult_out_1[108] + mult_out_2[108] + mult_out_3[108]) % 3329;
                                                                                                                                                                                 mul_add_t[2][109] <= (mult_out_1[109] + mult_out_2[109] + mult_out_3[109]) % 3329;
                                                                                                                                                                                 mul_add_t[2][110] <= (mult_out_1[110] + mult_out_2[110] + mult_out_3[110]) % 3329;
                                                                                                                                                                                 mul_add_t[2][111] <= (mult_out_1[111] + mult_out_2[111] + mult_out_3[111]) % 3329;
                                                                                                                                                                                 mul_add_t[2][112] <= (mult_out_1[112] + mult_out_2[112] + mult_out_3[112]) % 3329;
                                                                                                                                                                                 mul_add_t[2][113] <= (mult_out_1[113] + mult_out_2[113] + mult_out_3[113]) % 3329;
                                                                                                                                                                                 mul_add_t[2][114] <= (mult_out_1[114] + mult_out_2[114] + mult_out_3[114]) % 3329;
                                                                                                                                                                                 mul_add_t[2][115] <= (mult_out_1[115] + mult_out_2[115] + mult_out_3[115]) % 3329;
                                                                                                                                                                                 mul_add_t[2][116] <= (mult_out_1[116] + mult_out_2[116] + mult_out_3[116]) % 3329;
                                                                                                                                                                                 mul_add_t[2][117] <= (mult_out_1[117] + mult_out_2[117] + mult_out_3[117]) % 3329;
                                                                                                                                                                                 mul_add_t[2][118] <= (mult_out_1[118] + mult_out_2[118] + mult_out_3[118]) % 3329;
                                                                                                                                                                                 mul_add_t[2][119] <= (mult_out_1[119] + mult_out_2[119] + mult_out_3[119]) % 3329;
                                                                                                                                                                                 mul_add_t[2][120] <= (mult_out_1[120] + mult_out_2[120] + mult_out_3[120]) % 3329;
                                                                                                                                                                                 mul_add_t[2][121] <= (mult_out_1[121] + mult_out_2[121] + mult_out_3[121]) % 3329;
                                                                                                                                                                                 mul_add_t[2][122] <= (mult_out_1[122] + mult_out_2[122] + mult_out_3[122]) % 3329;
                                                                                                                                                                                 mul_add_t[2][123] <= (mult_out_1[123] + mult_out_2[123] + mult_out_3[123]) % 3329;
                                                                                                                                                                                 mul_add_t[2][124] <= (mult_out_1[124] + mult_out_2[124] + mult_out_3[124]) % 3329;
                                                                                                                                                                                 mul_add_t[2][125] <= (mult_out_1[125] + mult_out_2[125] + mult_out_3[125]) % 3329;
                                                                                                                                                                                 mul_add_t[2][126] <= (mult_out_1[126] + mult_out_2[126] + mult_out_3[126]) % 3329;
                                                                                                                                                                                 mul_add_t[2][127] <= (mult_out_1[127] + mult_out_2[127] + mult_out_3[127]) % 3329;
                                                                                                                                                                                 mul_add_t[2][128] <= (mult_out_1[128] + mult_out_2[128] + mult_out_3[128]) % 3329;
                                                                                                                                                                                 mul_add_t[2][129] <= (mult_out_1[129] + mult_out_2[129] + mult_out_3[129]) % 3329;
                                                                                                                                                                                 mul_add_t[2][130] <= (mult_out_1[130] + mult_out_2[130] + mult_out_3[130]) % 3329;
                                                                                                                                                                                 mul_add_t[2][131] <= (mult_out_1[131] + mult_out_2[131] + mult_out_3[131]) % 3329;
                                                                                                                                                                                 mul_add_t[2][132] <= (mult_out_1[132] + mult_out_2[132] + mult_out_3[132]) % 3329;
                                                                                                                                                                                 mul_add_t[2][133] <= (mult_out_1[133] + mult_out_2[133] + mult_out_3[133]) % 3329;
                                                                                                                                                                                 mul_add_t[2][134] <= (mult_out_1[134] + mult_out_2[134] + mult_out_3[134]) % 3329;
                                                                                                                                                                                 mul_add_t[2][135] <= (mult_out_1[135] + mult_out_2[135] + mult_out_3[135]) % 3329;
                                                                                                                                                                                 mul_add_t[2][136] <= (mult_out_1[136] + mult_out_2[136] + mult_out_3[136]) % 3329;
                                                                                                                                                                                 mul_add_t[2][137] <= (mult_out_1[137] + mult_out_2[137] + mult_out_3[137]) % 3329;
                                                                                                                                                                                 mul_add_t[2][138] <= (mult_out_1[138] + mult_out_2[138] + mult_out_3[138]) % 3329;
                                                                                                                                                                                 mul_add_t[2][139] <= (mult_out_1[139] + mult_out_2[139] + mult_out_3[139]) % 3329;
                                                                                                                                                                                 mul_add_t[2][140] <= (mult_out_1[140] + mult_out_2[140] + mult_out_3[140]) % 3329;
                                                                                                                                                                                 mul_add_t[2][141] <= (mult_out_1[141] + mult_out_2[141] + mult_out_3[141]) % 3329;
                                                                                                                                                                                 mul_add_t[2][142] <= (mult_out_1[142] + mult_out_2[142] + mult_out_3[142]) % 3329;
                                                                                                                                                                                 mul_add_t[2][143] <= (mult_out_1[143] + mult_out_2[143] + mult_out_3[143]) % 3329;
                                                                                                                                                                                 mul_add_t[2][144] <= (mult_out_1[144] + mult_out_2[144] + mult_out_3[144]) % 3329;
                                                                                                                                                                                 mul_add_t[2][145] <= (mult_out_1[145] + mult_out_2[145] + mult_out_3[145]) % 3329;
                                                                                                                                                                                 mul_add_t[2][146] <= (mult_out_1[146] + mult_out_2[146] + mult_out_3[146]) % 3329;
                                                                                                                                                                                 mul_add_t[2][147] <= (mult_out_1[147] + mult_out_2[147] + mult_out_3[147]) % 3329;
                                                                                                                                                                                 mul_add_t[2][148] <= (mult_out_1[148] + mult_out_2[148] + mult_out_3[148]) % 3329;
                                                                                                                                                                                 mul_add_t[2][149] <= (mult_out_1[149] + mult_out_2[149] + mult_out_3[149]) % 3329;
                                                                                                                                                                                 mul_add_t[2][150] <= (mult_out_1[150] + mult_out_2[150] + mult_out_3[150]) % 3329;
                                                                                                                                                                                 mul_add_t[2][151] <= (mult_out_1[151] + mult_out_2[151] + mult_out_3[151]) % 3329;
                                                                                                                                                                                 mul_add_t[2][152] <= (mult_out_1[152] + mult_out_2[152] + mult_out_3[152]) % 3329;
                                                                                                                                                                                 mul_add_t[2][153] <= (mult_out_1[153] + mult_out_2[153] + mult_out_3[153]) % 3329;
                                                                                                                                                                                 mul_add_t[2][154] <= (mult_out_1[154] + mult_out_2[154] + mult_out_3[154]) % 3329;
                                                                                                                                                                                 mul_add_t[2][155] <= (mult_out_1[155] + mult_out_2[155] + mult_out_3[155]) % 3329;
                                                                                                                                                                                 mul_add_t[2][156] <= (mult_out_1[156] + mult_out_2[156] + mult_out_3[156]) % 3329;
                                                                                                                                                                                 mul_add_t[2][157] <= (mult_out_1[157] + mult_out_2[157] + mult_out_3[157]) % 3329;
                                                                                                                                                                                 mul_add_t[2][158] <= (mult_out_1[158] + mult_out_2[158] + mult_out_3[158]) % 3329;
                                                                                                                                                                                 mul_add_t[2][159] <= (mult_out_1[159] + mult_out_2[159] + mult_out_3[159]) % 3329;
                                                                                                                                                                                 mul_add_t[2][160] <= (mult_out_1[160] + mult_out_2[160] + mult_out_3[160]) % 3329;
                                                                                                                                                                                 mul_add_t[2][161] <= (mult_out_1[161] + mult_out_2[161] + mult_out_3[161]) % 3329;
                                                                                                                                                                                 mul_add_t[2][162] <= (mult_out_1[162] + mult_out_2[162] + mult_out_3[162]) % 3329;
                                                                                                                                                                                 mul_add_t[2][163] <= (mult_out_1[163] + mult_out_2[163] + mult_out_3[163]) % 3329;
                                                                                                                                                                                 mul_add_t[2][164] <= (mult_out_1[164] + mult_out_2[164] + mult_out_3[164]) % 3329;
                                                                                                                                                                                 mul_add_t[2][165] <= (mult_out_1[165] + mult_out_2[165] + mult_out_3[165]) % 3329;
                                                                                                                                                                                 mul_add_t[2][166] <= (mult_out_1[166] + mult_out_2[166] + mult_out_3[166]) % 3329;
                                                                                                                                                                                 mul_add_t[2][167] <= (mult_out_1[167] + mult_out_2[167] + mult_out_3[167]) % 3329;
                                                                                                                                                                                 mul_add_t[2][168] <= (mult_out_1[168] + mult_out_2[168] + mult_out_3[168]) % 3329;
                                                                                                                                                                                 mul_add_t[2][169] <= (mult_out_1[169] + mult_out_2[169] + mult_out_3[169]) % 3329;
                                                                                                                                                                                 mul_add_t[2][170] <= (mult_out_1[170] + mult_out_2[170] + mult_out_3[170]) % 3329;
                                                                                                                                                                                 mul_add_t[2][171] <= (mult_out_1[171] + mult_out_2[171] + mult_out_3[171]) % 3329;
                                                                                                                                                                                 mul_add_t[2][172] <= (mult_out_1[172] + mult_out_2[172] + mult_out_3[172]) % 3329;
                                                                                                                                                                                 mul_add_t[2][173] <= (mult_out_1[173] + mult_out_2[173] + mult_out_3[173]) % 3329;
                                                                                                                                                                                 mul_add_t[2][174] <= (mult_out_1[174] + mult_out_2[174] + mult_out_3[174]) % 3329;
                                                                                                                                                                                 mul_add_t[2][175] <= (mult_out_1[175] + mult_out_2[175] + mult_out_3[175]) % 3329;
                                                                                                                                                                                 mul_add_t[2][176] <= (mult_out_1[176] + mult_out_2[176] + mult_out_3[176]) % 3329;
                                                                                                                                                                                 mul_add_t[2][177] <= (mult_out_1[177] + mult_out_2[177] + mult_out_3[177]) % 3329;
                                                                                                                                                                                 mul_add_t[2][178] <= (mult_out_1[178] + mult_out_2[178] + mult_out_3[178]) % 3329;
                                                                                                                                                                                 mul_add_t[2][179] <= (mult_out_1[179] + mult_out_2[179] + mult_out_3[179]) % 3329;
                                                                                                                                                                                 mul_add_t[2][180] <= (mult_out_1[180] + mult_out_2[180] + mult_out_3[180]) % 3329;
                                                                                                                                                                                 mul_add_t[2][181] <= (mult_out_1[181] + mult_out_2[181] + mult_out_3[181]) % 3329;
                                                                                                                                                                                 mul_add_t[2][182] <= (mult_out_1[182] + mult_out_2[182] + mult_out_3[182]) % 3329;
                                                                                                                                                                                 mul_add_t[2][183] <= (mult_out_1[183] + mult_out_2[183] + mult_out_3[183]) % 3329;
                                                                                                                                                                                 mul_add_t[2][184] <= (mult_out_1[184] + mult_out_2[184] + mult_out_3[184]) % 3329;
                                                                                                                                                                                 mul_add_t[2][185] <= (mult_out_1[185] + mult_out_2[185] + mult_out_3[185]) % 3329;
                                                                                                                                                                                 mul_add_t[2][186] <= (mult_out_1[186] + mult_out_2[186] + mult_out_3[186]) % 3329;
                                                                                                                                                                                 mul_add_t[2][187] <= (mult_out_1[187] + mult_out_2[187] + mult_out_3[187]) % 3329;
                                                                                                                                                                                 mul_add_t[2][188] <= (mult_out_1[188] + mult_out_2[188] + mult_out_3[188]) % 3329;
                                                                                                                                                                                 mul_add_t[2][189] <= (mult_out_1[189] + mult_out_2[189] + mult_out_3[189]) % 3329;
                                                                                                                                                                                 mul_add_t[2][190] <= (mult_out_1[190] + mult_out_2[190] + mult_out_3[190]) % 3329;
                                                                                                                                                                                 mul_add_t[2][191] <= (mult_out_1[191] + mult_out_2[191] + mult_out_3[191]) % 3329;
                                                                                                                                                                                 mul_add_t[2][192] <= (mult_out_1[192] + mult_out_2[192] + mult_out_3[192]) % 3329;
                                                                                                                                                                                 mul_add_t[2][193] <= (mult_out_1[193] + mult_out_2[193] + mult_out_3[193]) % 3329;
                                                                                                                                                                                 mul_add_t[2][194] <= (mult_out_1[194] + mult_out_2[194] + mult_out_3[194]) % 3329;
                                                                                                                                                                                 mul_add_t[2][195] <= (mult_out_1[195] + mult_out_2[195] + mult_out_3[195]) % 3329;
                                                                                                                                                                                 mul_add_t[2][196] <= (mult_out_1[196] + mult_out_2[196] + mult_out_3[196]) % 3329;
                                                                                                                                                                                 mul_add_t[2][197] <= (mult_out_1[197] + mult_out_2[197] + mult_out_3[197]) % 3329;
                                                                                                                                                                                 mul_add_t[2][198] <= (mult_out_1[198] + mult_out_2[198] + mult_out_3[198]) % 3329;
                                                                                                                                                                                 mul_add_t[2][199] <= (mult_out_1[199] + mult_out_2[199] + mult_out_3[199]) % 3329;
                                                                                                                                                                                 mul_add_t[2][200] <= (mult_out_1[200] + mult_out_2[200] + mult_out_3[200]) % 3329;
                                                                                                                                                                                 mul_add_t[2][201] <= (mult_out_1[201] + mult_out_2[201] + mult_out_3[201]) % 3329;
                                                                                                                                                                                 mul_add_t[2][202] <= (mult_out_1[202] + mult_out_2[202] + mult_out_3[202]) % 3329;
                                                                                                                                                                                 mul_add_t[2][203] <= (mult_out_1[203] + mult_out_2[203] + mult_out_3[203]) % 3329;
                                                                                                                                                                                 mul_add_t[2][204] <= (mult_out_1[204] + mult_out_2[204] + mult_out_3[204]) % 3329;
                                                                                                                                                                                 mul_add_t[2][205] <= (mult_out_1[205] + mult_out_2[205] + mult_out_3[205]) % 3329;
                                                                                                                                                                                 mul_add_t[2][206] <= (mult_out_1[206] + mult_out_2[206] + mult_out_3[206]) % 3329;
                                                                                                                                                                                 mul_add_t[2][207] <= (mult_out_1[207] + mult_out_2[207] + mult_out_3[207]) % 3329;
                                                                                                                                                                                 mul_add_t[2][208] <= (mult_out_1[208] + mult_out_2[208] + mult_out_3[208]) % 3329;
                                                                                                                                                                                 mul_add_t[2][209] <= (mult_out_1[209] + mult_out_2[209] + mult_out_3[209]) % 3329;
                                                                                                                                                                                 mul_add_t[2][210] <= (mult_out_1[210] + mult_out_2[210] + mult_out_3[210]) % 3329;
                                                                                                                                                                                 mul_add_t[2][211] <= (mult_out_1[211] + mult_out_2[211] + mult_out_3[211]) % 3329;
                                                                                                                                                                                 mul_add_t[2][212] <= (mult_out_1[212] + mult_out_2[212] + mult_out_3[212]) % 3329;
                                                                                                                                                                                 mul_add_t[2][213] <= (mult_out_1[213] + mult_out_2[213] + mult_out_3[213]) % 3329;
                                                                                                                                                                                 mul_add_t[2][214] <= (mult_out_1[214] + mult_out_2[214] + mult_out_3[214]) % 3329;
                                                                                                                                                                                 mul_add_t[2][215] <= (mult_out_1[215] + mult_out_2[215] + mult_out_3[215]) % 3329;
                                                                                                                                                                                 mul_add_t[2][216] <= (mult_out_1[216] + mult_out_2[216] + mult_out_3[216]) % 3329;
                                                                                                                                                                                 mul_add_t[2][217] <= (mult_out_1[217] + mult_out_2[217] + mult_out_3[217]) % 3329;
                                                                                                                                                                                 mul_add_t[2][218] <= (mult_out_1[218] + mult_out_2[218] + mult_out_3[218]) % 3329;
                                                                                                                                                                                 mul_add_t[2][219] <= (mult_out_1[219] + mult_out_2[219] + mult_out_3[219]) % 3329;
                                                                                                                                                                                 mul_add_t[2][220] <= (mult_out_1[220] + mult_out_2[220] + mult_out_3[220]) % 3329;
                                                                                                                                                                                 mul_add_t[2][221] <= (mult_out_1[221] + mult_out_2[221] + mult_out_3[221]) % 3329;
                                                                                                                                                                                 mul_add_t[2][222] <= (mult_out_1[222] + mult_out_2[222] + mult_out_3[222]) % 3329;
                                                                                                                                                                                 mul_add_t[2][223] <= (mult_out_1[223] + mult_out_2[223] + mult_out_3[223]) % 3329;
                                                                                                                                                                                 mul_add_t[2][224] <= (mult_out_1[224] + mult_out_2[224] + mult_out_3[224]) % 3329;
                                                                                                                                                                                 mul_add_t[2][225] <= (mult_out_1[225] + mult_out_2[225] + mult_out_3[225]) % 3329;
                                                                                                                                                                                 mul_add_t[2][226] <= (mult_out_1[226] + mult_out_2[226] + mult_out_3[226]) % 3329;
                                                                                                                                                                                 mul_add_t[2][227] <= (mult_out_1[227] + mult_out_2[227] + mult_out_3[227]) % 3329;
                                                                                                                                                                                 mul_add_t[2][228] <= (mult_out_1[228] + mult_out_2[228] + mult_out_3[228]) % 3329;
                                                                                                                                                                                 mul_add_t[2][229] <= (mult_out_1[229] + mult_out_2[229] + mult_out_3[229]) % 3329;
                                                                                                                                                                                 mul_add_t[2][230] <= (mult_out_1[230] + mult_out_2[230] + mult_out_3[230]) % 3329;
                                                                                                                                                                                 mul_add_t[2][231] <= (mult_out_1[231] + mult_out_2[231] + mult_out_3[231]) % 3329;
                                                                                                                                                                                 mul_add_t[2][232] <= (mult_out_1[232] + mult_out_2[232] + mult_out_3[232]) % 3329;
                                                                                                                                                                                 mul_add_t[2][233] <= (mult_out_1[233] + mult_out_2[233] + mult_out_3[233]) % 3329;
                                                                                                                                                                                 mul_add_t[2][234] <= (mult_out_1[234] + mult_out_2[234] + mult_out_3[234]) % 3329;
                                                                                                                                                                                 mul_add_t[2][235] <= (mult_out_1[235] + mult_out_2[235] + mult_out_3[235]) % 3329;
                                                                                                                                                                                 mul_add_t[2][236] <= (mult_out_1[236] + mult_out_2[236] + mult_out_3[236]) % 3329;
                                                                                                                                                                                 mul_add_t[2][237] <= (mult_out_1[237] + mult_out_2[237] + mult_out_3[237]) % 3329;
                                                                                                                                                                                 mul_add_t[2][238] <= (mult_out_1[238] + mult_out_2[238] + mult_out_3[238]) % 3329;
                                                                                                                                                                                 mul_add_t[2][239] <= (mult_out_1[239] + mult_out_2[239] + mult_out_3[239]) % 3329;
                                                                                                                                                                                 mul_add_t[2][240] <= (mult_out_1[240] + mult_out_2[240] + mult_out_3[240]) % 3329;
                                                                                                                                                                                 mul_add_t[2][241] <= (mult_out_1[241] + mult_out_2[241] + mult_out_3[241]) % 3329;
                                                                                                                                                                                 mul_add_t[2][242] <= (mult_out_1[242] + mult_out_2[242] + mult_out_3[242]) % 3329;
                                                                                                                                                                                 mul_add_t[2][243] <= (mult_out_1[243] + mult_out_2[243] + mult_out_3[243]) % 3329;
                                                                                                                                                                                 mul_add_t[2][244] <= (mult_out_1[244] + mult_out_2[244] + mult_out_3[244]) % 3329;
                                                                                                                                                                                 mul_add_t[2][245] <= (mult_out_1[245] + mult_out_2[245] + mult_out_3[245]) % 3329;
                                                                                                                                                                                 mul_add_t[2][246] <= (mult_out_1[246] + mult_out_2[246] + mult_out_3[246]) % 3329;
                                                                                                                                                                                 mul_add_t[2][247] <= (mult_out_1[247] + mult_out_2[247] + mult_out_3[247]) % 3329;
                                                                                                                                                                                 mul_add_t[2][248] <= (mult_out_1[248] + mult_out_2[248] + mult_out_3[248]) % 3329;
                                                                                                                                                                                 mul_add_t[2][249] <= (mult_out_1[249] + mult_out_2[249] + mult_out_3[249]) % 3329;
                                                                                                                                                                                 mul_add_t[2][250] <= (mult_out_1[250] + mult_out_2[250] + mult_out_3[250]) % 3329;
                                                                                                                                                                                 mul_add_t[2][251] <= (mult_out_1[251] + mult_out_2[251] + mult_out_3[251]) % 3329;
                                                                                                                                                                                 mul_add_t[2][252] <= (mult_out_1[252] + mult_out_2[252] + mult_out_3[252]) % 3329;
                                                                                                                                                                                 mul_add_t[2][253] <= (mult_out_1[253] + mult_out_2[253] + mult_out_3[253]) % 3329;
                                                                                                                                                                                 mul_add_t[2][254] <= (mult_out_1[254] + mult_out_2[254] + mult_out_3[254]) % 3329;
                                                                                                                                                                                 mul_add_t[2][255] <= (mult_out_1[255] + mult_out_2[255] + mult_out_3[255]) % 3329;
                                                                                                                                                                                 u[0][0] = in_1[0] + e1[0][0] %3329;
                                                                                                                                                                                 u[0][1] = in_1[1] + e1[0][1] %3329;
                                                                                                                                                                                 u[0][2] = in_1[2] + e1[0][2] %3329;
                                                                                                                                                                                 u[0][3] = in_1[3] + e1[0][3] %3329;
                                                                                                                                                                                 u[0][4] = in_1[4] + e1[0][4] %3329;
                                                                                                                                                                                 u[0][5] = in_1[5] + e1[0][5] %3329;
                                                                                                                                                                                 u[0][6] = in_1[6] + e1[0][6] %3329;
                                                                                                                                                                                 u[0][7] = in_1[7] + e1[0][7] %3329;
                                                                                                                                                                                 u[0][8] = in_1[8] + e1[0][8] %3329;
                                                                                                                                                                                 u[0][9] = in_1[9] + e1[0][9] %3329;
                                                                                                                                                                                 u[0][10] = in_1[10] + e1[0][10] %3329;
                                                                                                                                                                                 u[0][11] = in_1[11] + e1[0][11] %3329;
                                                                                                                                                                                 u[0][12] = in_1[12] + e1[0][12] %3329;
                                                                                                                                                                                 u[0][13] = in_1[13] + e1[0][13] %3329;
                                                                                                                                                                                 u[0][14] = in_1[14] + e1[0][14] %3329;
                                                                                                                                                                                 u[0][15] = in_1[15] + e1[0][15] %3329;
                                                                                                                                                                                 u[0][16] = in_1[16] + e1[0][16] %3329;
                                                                                                                                                                                 u[0][17] = in_1[17] + e1[0][17] %3329;
                                                                                                                                                                                 u[0][18] = in_1[18] + e1[0][18] %3329;
                                                                                                                                                                                 u[0][19] = in_1[19] + e1[0][19] %3329;
                                                                                                                                                                                 u[0][20] = in_1[20] + e1[0][20] %3329;
                                                                                                                                                                                 u[0][21] = in_1[21] + e1[0][21] %3329;
                                                                                                                                                                                 u[0][22] = in_1[22] + e1[0][22] %3329;
                                                                                                                                                                                 u[0][23] = in_1[23] + e1[0][23] %3329;
                                                                                                                                                                                 u[0][24] = in_1[24] + e1[0][24] %3329;
                                                                                                                                                                                 u[0][25] = in_1[25] + e1[0][25] %3329;
                                                                                                                                                                                 u[0][26] = in_1[26] + e1[0][26] %3329;
                                                                                                                                                                                 u[0][27] = in_1[27] + e1[0][27] %3329;
                                                                                                                                                                                 u[0][28] = in_1[28] + e1[0][28] %3329;
                                                                                                                                                                                 u[0][29] = in_1[29] + e1[0][29] %3329;
                                                                                                                                                                                 u[0][30] = in_1[30] + e1[0][30] %3329;
                                                                                                                                                                                 u[0][31] = in_1[31] + e1[0][31] %3329;
                                                                                                                                                                                 u[0][32] = in_1[32] + e1[0][32] %3329;
                                                                                                                                                                                 u[0][33] = in_1[33] + e1[0][33] %3329;
                                                                                                                                                                                 u[0][34] = in_1[34] + e1[0][34] %3329;
                                                                                                                                                                                 u[0][35] = in_1[35] + e1[0][35] %3329;
                                                                                                                                                                                 u[0][36] = in_1[36] + e1[0][36] %3329;
                                                                                                                                                                                 u[0][37] = in_1[37] + e1[0][37] %3329;
                                                                                                                                                                                 u[0][38] = in_1[38] + e1[0][38] %3329;
                                                                                                                                                                                 u[0][39] = in_1[39] + e1[0][39] %3329;
                                                                                                                                                                                 u[0][40] = in_1[40] + e1[0][40] %3329;
                                                                                                                                                                                 u[0][41] = in_1[41] + e1[0][41] %3329;
                                                                                                                                                                                 u[0][42] = in_1[42] + e1[0][42] %3329;
                                                                                                                                                                                 u[0][43] = in_1[43] + e1[0][43] %3329;
                                                                                                                                                                                 u[0][44] = in_1[44] + e1[0][44] %3329;
                                                                                                                                                                                 u[0][45] = in_1[45] + e1[0][45] %3329;
                                                                                                                                                                                 u[0][46] = in_1[46] + e1[0][46] %3329;
                                                                                                                                                                                 u[0][47] = in_1[47] + e1[0][47] %3329;
                                                                                                                                                                                 u[0][48] = in_1[48] + e1[0][48] %3329;
                                                                                                                                                                                 u[0][49] = in_1[49] + e1[0][49] %3329;
                                                                                                                                                                                 u[0][50] = in_1[50] + e1[0][50] %3329;
                                                                                                                                                                                 u[0][51] = in_1[51] + e1[0][51] %3329;
                                                                                                                                                                                 u[0][52] = in_1[52] + e1[0][52] %3329;
                                                                                                                                                                                 u[0][53] = in_1[53] + e1[0][53] %3329;
                                                                                                                                                                                 u[0][54] = in_1[54] + e1[0][54] %3329;
                                                                                                                                                                                 u[0][55] = in_1[55] + e1[0][55] %3329;
                                                                                                                                                                                 u[0][56] = in_1[56] + e1[0][56] %3329;
                                                                                                                                                                                 u[0][57] = in_1[57] + e1[0][57] %3329;
                                                                                                                                                                                 u[0][58] = in_1[58] + e1[0][58] %3329;
                                                                                                                                                                                 u[0][59] = in_1[59] + e1[0][59] %3329;
                                                                                                                                                                                 u[0][60] = in_1[60] + e1[0][60] %3329;
                                                                                                                                                                                 u[0][61] = in_1[61] + e1[0][61] %3329;
                                                                                                                                                                                 u[0][62] = in_1[62] + e1[0][62] %3329;
                                                                                                                                                                                 u[0][63] = in_1[63] + e1[0][63] %3329;
                                                                                                                                                                                 u[0][64] = in_1[64] + e1[0][64] %3329;
                                                                                                                                                                                 u[0][65] = in_1[65] + e1[0][65] %3329;
                                                                                                                                                                                 u[0][66] = in_1[66] + e1[0][66] %3329;
                                                                                                                                                                                 u[0][67] = in_1[67] + e1[0][67] %3329;
                                                                                                                                                                                 u[0][68] = in_1[68] + e1[0][68] %3329;
                                                                                                                                                                                 u[0][69] = in_1[69] + e1[0][69] %3329;
                                                                                                                                                                                 u[0][70] = in_1[70] + e1[0][70] %3329;
                                                                                                                                                                                 u[0][71] = in_1[71] + e1[0][71] %3329;
                                                                                                                                                                                 u[0][72] = in_1[72] + e1[0][72] %3329;
                                                                                                                                                                                 u[0][73] = in_1[73] + e1[0][73] %3329;
                                                                                                                                                                                 u[0][74] = in_1[74] + e1[0][74] %3329;
                                                                                                                                                                                 u[0][75] = in_1[75] + e1[0][75] %3329;
                                                                                                                                                                                 u[0][76] = in_1[76] + e1[0][76] %3329;
                                                                                                                                                                                 u[0][77] = in_1[77] + e1[0][77] %3329;
                                                                                                                                                                                 u[0][78] = in_1[78] + e1[0][78] %3329;
                                                                                                                                                                                 u[0][79] = in_1[79] + e1[0][79] %3329;
                                                                                                                                                                                 u[0][80] = in_1[80] + e1[0][80] %3329;
                                                                                                                                                                                 u[0][81] = in_1[81] + e1[0][81] %3329;
                                                                                                                                                                                 u[0][82] = in_1[82] + e1[0][82] %3329;
                                                                                                                                                                                 u[0][83] = in_1[83] + e1[0][83] %3329;
                                                                                                                                                                                 u[0][84] = in_1[84] + e1[0][84] %3329;
                                                                                                                                                                                 u[0][85] = in_1[85] + e1[0][85] %3329;
                                                                                                                                                                                 u[0][86] = in_1[86] + e1[0][86] %3329;
                                                                                                                                                                                 u[0][87] = in_1[87] + e1[0][87] %3329;
                                                                                                                                                                                 u[0][88] = in_1[88] + e1[0][88] %3329;
                                                                                                                                                                                 u[0][89] = in_1[89] + e1[0][89] %3329;
                                                                                                                                                                                 u[0][90] = in_1[90] + e1[0][90] %3329;
                                                                                                                                                                                 u[0][91] = in_1[91] + e1[0][91] %3329;
                                                                                                                                                                                 u[0][92] = in_1[92] + e1[0][92] %3329;
                                                                                                                                                                                 u[0][93] = in_1[93] + e1[0][93] %3329;
                                                                                                                                                                                 u[0][94] = in_1[94] + e1[0][94] %3329;
                                                                                                                                                                                 u[0][95] = in_1[95] + e1[0][95] %3329;
                                                                                                                                                                                 u[0][96] = in_1[96] + e1[0][96] %3329;
                                                                                                                                                                                 u[0][97] = in_1[97] + e1[0][97] %3329;
                                                                                                                                                                                 u[0][98] = in_1[98] + e1[0][98] %3329;
                                                                                                                                                                                 u[0][99] = in_1[99] + e1[0][99] %3329;
                                                                                                                                                                                 u[0][100] = in_1[100] + e1[0][100] %3329;
                                                                                                                                                                                 u[0][101] = in_1[101] + e1[0][101] %3329;
                                                                                                                                                                                 u[0][102] = in_1[102] + e1[0][102] %3329;
                                                                                                                                                                                 u[0][103] = in_1[103] + e1[0][103] %3329;
                                                                                                                                                                                 u[0][104] = in_1[104] + e1[0][104] %3329;
                                                                                                                                                                                 u[0][105] = in_1[105] + e1[0][105] %3329;
                                                                                                                                                                                 u[0][106] = in_1[106] + e1[0][106] %3329;
                                                                                                                                                                                 u[0][107] = in_1[107] + e1[0][107] %3329;
                                                                                                                                                                                 u[0][108] = in_1[108] + e1[0][108] %3329;
                                                                                                                                                                                 u[0][109] = in_1[109] + e1[0][109] %3329;
                                                                                                                                                                                 u[0][110] = in_1[110] + e1[0][110] %3329;
                                                                                                                                                                                 u[0][111] = in_1[111] + e1[0][111] %3329;
                                                                                                                                                                                 u[0][112] = in_1[112] + e1[0][112] %3329;
                                                                                                                                                                                 u[0][113] = in_1[113] + e1[0][113] %3329;
                                                                                                                                                                                 u[0][114] = in_1[114] + e1[0][114] %3329;
                                                                                                                                                                                 u[0][115] = in_1[115] + e1[0][115] %3329;
                                                                                                                                                                                 u[0][116] = in_1[116] + e1[0][116] %3329;
                                                                                                                                                                                 u[0][117] = in_1[117] + e1[0][117] %3329;
                                                                                                                                                                                 u[0][118] = in_1[118] + e1[0][118] %3329;
                                                                                                                                                                                 u[0][119] = in_1[119] + e1[0][119] %3329;
                                                                                                                                                                                 u[0][120] = in_1[120] + e1[0][120] %3329;
                                                                                                                                                                                 u[0][121] = in_1[121] + e1[0][121] %3329;
                                                                                                                                                                                 u[0][122] = in_1[122] + e1[0][122] %3329;
                                                                                                                                                                                 u[0][123] = in_1[123] + e1[0][123] %3329;
                                                                                                                                                                                 u[0][124] = in_1[124] + e1[0][124] %3329;
                                                                                                                                                                                 u[0][125] = in_1[125] + e1[0][125] %3329;
                                                                                                                                                                                 u[0][126] = in_1[126] + e1[0][126] %3329;
                                                                                                                                                                                 u[0][127] = in_1[127] + e1[0][127] %3329;
                                                                                                                                                                                 u[0][128] = in_1[128] + e1[0][128] %3329;
                                                                                                                                                                                 u[0][129] = in_1[129] + e1[0][129] %3329;
                                                                                                                                                                                 u[0][130] = in_1[130] + e1[0][130] %3329;
                                                                                                                                                                                 u[0][131] = in_1[131] + e1[0][131] %3329;
                                                                                                                                                                                 u[0][132] = in_1[132] + e1[0][132] %3329;
                                                                                                                                                                                 u[0][133] = in_1[133] + e1[0][133] %3329;
                                                                                                                                                                                 u[0][134] = in_1[134] + e1[0][134] %3329;
                                                                                                                                                                                 u[0][135] = in_1[135] + e1[0][135] %3329;
                                                                                                                                                                                 u[0][136] = in_1[136] + e1[0][136] %3329;
                                                                                                                                                                                 u[0][137] = in_1[137] + e1[0][137] %3329;
                                                                                                                                                                                 u[0][138] = in_1[138] + e1[0][138] %3329;
                                                                                                                                                                                 u[0][139] = in_1[139] + e1[0][139] %3329;
                                                                                                                                                                                 u[0][140] = in_1[140] + e1[0][140] %3329;
                                                                                                                                                                                 u[0][141] = in_1[141] + e1[0][141] %3329;
                                                                                                                                                                                 u[0][142] = in_1[142] + e1[0][142] %3329;
                                                                                                                                                                                 u[0][143] = in_1[143] + e1[0][143] %3329;
                                                                                                                                                                                 u[0][144] = in_1[144] + e1[0][144] %3329;
                                                                                                                                                                                 u[0][145] = in_1[145] + e1[0][145] %3329;
                                                                                                                                                                                 u[0][146] = in_1[146] + e1[0][146] %3329;
                                                                                                                                                                                 u[0][147] = in_1[147] + e1[0][147] %3329;
                                                                                                                                                                                 u[0][148] = in_1[148] + e1[0][148] %3329;
                                                                                                                                                                                 u[0][149] = in_1[149] + e1[0][149] %3329;
                                                                                                                                                                                 u[0][150] = in_1[150] + e1[0][150] %3329;
                                                                                                                                                                                 u[0][151] = in_1[151] + e1[0][151] %3329;
                                                                                                                                                                                 u[0][152] = in_1[152] + e1[0][152] %3329;
                                                                                                                                                                                 u[0][153] = in_1[153] + e1[0][153] %3329;
                                                                                                                                                                                 u[0][154] = in_1[154] + e1[0][154] %3329;
                                                                                                                                                                                 u[0][155] = in_1[155] + e1[0][155] %3329;
                                                                                                                                                                                 u[0][156] = in_1[156] + e1[0][156] %3329;
                                                                                                                                                                                 u[0][157] = in_1[157] + e1[0][157] %3329;
                                                                                                                                                                                 u[0][158] = in_1[158] + e1[0][158] %3329;
                                                                                                                                                                                 u[0][159] = in_1[159] + e1[0][159] %3329;
                                                                                                                                                                                 u[0][160] = in_1[160] + e1[0][160] %3329;
                                                                                                                                                                                 u[0][161] = in_1[161] + e1[0][161] %3329;
                                                                                                                                                                                 u[0][162] = in_1[162] + e1[0][162] %3329;
                                                                                                                                                                                 u[0][163] = in_1[163] + e1[0][163] %3329;
                                                                                                                                                                                 u[0][164] = in_1[164] + e1[0][164] %3329;
                                                                                                                                                                                 u[0][165] = in_1[165] + e1[0][165] %3329;
                                                                                                                                                                                 u[0][166] = in_1[166] + e1[0][166] %3329;
                                                                                                                                                                                 u[0][167] = in_1[167] + e1[0][167] %3329;
                                                                                                                                                                                 u[0][168] = in_1[168] + e1[0][168] %3329;
                                                                                                                                                                                 u[0][169] = in_1[169] + e1[0][169] %3329;
                                                                                                                                                                                 u[0][170] = in_1[170] + e1[0][170] %3329;
                                                                                                                                                                                 u[0][171] = in_1[171] + e1[0][171] %3329;
                                                                                                                                                                                 u[0][172] = in_1[172] + e1[0][172] %3329;
                                                                                                                                                                                 u[0][173] = in_1[173] + e1[0][173] %3329;
                                                                                                                                                                                 u[0][174] = in_1[174] + e1[0][174] %3329;
                                                                                                                                                                                 u[0][175] = in_1[175] + e1[0][175] %3329;
                                                                                                                                                                                 u[0][176] = in_1[176] + e1[0][176] %3329;
                                                                                                                                                                                 u[0][177] = in_1[177] + e1[0][177] %3329;
                                                                                                                                                                                 u[0][178] = in_1[178] + e1[0][178] %3329;
                                                                                                                                                                                 u[0][179] = in_1[179] + e1[0][179] %3329;
                                                                                                                                                                                 u[0][180] = in_1[180] + e1[0][180] %3329;
                                                                                                                                                                                 u[0][181] = in_1[181] + e1[0][181] %3329;
                                                                                                                                                                                 u[0][182] = in_1[182] + e1[0][182] %3329;
                                                                                                                                                                                 u[0][183] = in_1[183] + e1[0][183] %3329;
                                                                                                                                                                                 u[0][184] = in_1[184] + e1[0][184] %3329;
                                                                                                                                                                                 u[0][185] = in_1[185] + e1[0][185] %3329;
                                                                                                                                                                                 u[0][186] = in_1[186] + e1[0][186] %3329;
                                                                                                                                                                                 u[0][187] = in_1[187] + e1[0][187] %3329;
                                                                                                                                                                                 u[0][188] = in_1[188] + e1[0][188] %3329;
                                                                                                                                                                                 u[0][189] = in_1[189] + e1[0][189] %3329;
                                                                                                                                                                                 u[0][190] = in_1[190] + e1[0][190] %3329;
                                                                                                                                                                                 u[0][191] = in_1[191] + e1[0][191] %3329;
                                                                                                                                                                                 u[0][192] = in_1[192] + e1[0][192] %3329;
                                                                                                                                                                                 u[0][193] = in_1[193] + e1[0][193] %3329;
                                                                                                                                                                                 u[0][194] = in_1[194] + e1[0][194] %3329;
                                                                                                                                                                                 u[0][195] = in_1[195] + e1[0][195] %3329;
                                                                                                                                                                                 u[0][196] = in_1[196] + e1[0][196] %3329;
                                                                                                                                                                                 u[0][197] = in_1[197] + e1[0][197] %3329;
                                                                                                                                                                                 u[0][198] = in_1[198] + e1[0][198] %3329;
                                                                                                                                                                                 u[0][199] = in_1[199] + e1[0][199] %3329;
                                                                                                                                                                                 u[0][200] = in_1[200] + e1[0][200] %3329;
                                                                                                                                                                                 u[0][201] = in_1[201] + e1[0][201] %3329;
                                                                                                                                                                                 u[0][202] = in_1[202] + e1[0][202] %3329;
                                                                                                                                                                                 u[0][203] = in_1[203] + e1[0][203] %3329;
                                                                                                                                                                                 u[0][204] = in_1[204] + e1[0][204] %3329;
                                                                                                                                                                                 u[0][205] = in_1[205] + e1[0][205] %3329;
                                                                                                                                                                                 u[0][206] = in_1[206] + e1[0][206] %3329;
                                                                                                                                                                                 u[0][207] = in_1[207] + e1[0][207] %3329;
                                                                                                                                                                                 u[0][208] = in_1[208] + e1[0][208] %3329;
                                                                                                                                                                                 u[0][209] = in_1[209] + e1[0][209] %3329;
                                                                                                                                                                                 u[0][210] = in_1[210] + e1[0][210] %3329;
                                                                                                                                                                                 u[0][211] = in_1[211] + e1[0][211] %3329;
                                                                                                                                                                                 u[0][212] = in_1[212] + e1[0][212] %3329;
                                                                                                                                                                                 u[0][213] = in_1[213] + e1[0][213] %3329;
                                                                                                                                                                                 u[0][214] = in_1[214] + e1[0][214] %3329;
                                                                                                                                                                                 u[0][215] = in_1[215] + e1[0][215] %3329;
                                                                                                                                                                                 u[0][216] = in_1[216] + e1[0][216] %3329;
                                                                                                                                                                                 u[0][217] = in_1[217] + e1[0][217] %3329;
                                                                                                                                                                                 u[0][218] = in_1[218] + e1[0][218] %3329;
                                                                                                                                                                                 u[0][219] = in_1[219] + e1[0][219] %3329;
                                                                                                                                                                                 u[0][220] = in_1[220] + e1[0][220] %3329;
                                                                                                                                                                                 u[0][221] = in_1[221] + e1[0][221] %3329;
                                                                                                                                                                                 u[0][222] = in_1[222] + e1[0][222] %3329;
                                                                                                                                                                                 u[0][223] = in_1[223] + e1[0][223] %3329;
                                                                                                                                                                                 u[0][224] = in_1[224] + e1[0][224] %3329;
                                                                                                                                                                                 u[0][225] = in_1[225] + e1[0][225] %3329;
                                                                                                                                                                                 u[0][226] = in_1[226] + e1[0][226] %3329;
                                                                                                                                                                                 u[0][227] = in_1[227] + e1[0][227] %3329;
                                                                                                                                                                                 u[0][228] = in_1[228] + e1[0][228] %3329;
                                                                                                                                                                                 u[0][229] = in_1[229] + e1[0][229] %3329;
                                                                                                                                                                                 u[0][230] = in_1[230] + e1[0][230] %3329;
                                                                                                                                                                                 u[0][231] = in_1[231] + e1[0][231] %3329;
                                                                                                                                                                                 u[0][232] = in_1[232] + e1[0][232] %3329;
                                                                                                                                                                                 u[0][233] = in_1[233] + e1[0][233] %3329;
                                                                                                                                                                                 u[0][234] = in_1[234] + e1[0][234] %3329;
                                                                                                                                                                                 u[0][235] = in_1[235] + e1[0][235] %3329;
                                                                                                                                                                                 u[0][236] = in_1[236] + e1[0][236] %3329;
                                                                                                                                                                                 u[0][237] = in_1[237] + e1[0][237] %3329;
                                                                                                                                                                                 u[0][238] = in_1[238] + e1[0][238] %3329;
                                                                                                                                                                                 u[0][239] = in_1[239] + e1[0][239] %3329;
                                                                                                                                                                                 u[0][240] = in_1[240] + e1[0][240] %3329;
                                                                                                                                                                                 u[0][241] = in_1[241] + e1[0][241] %3329;
                                                                                                                                                                                 u[0][242] = in_1[242] + e1[0][242] %3329;
                                                                                                                                                                                 u[0][243] = in_1[243] + e1[0][243] %3329;
                                                                                                                                                                                 u[0][244] = in_1[244] + e1[0][244] %3329;
                                                                                                                                                                                 u[0][245] = in_1[245] + e1[0][245] %3329;
                                                                                                                                                                                 u[0][246] = in_1[246] + e1[0][246] %3329;
                                                                                                                                                                                 u[0][247] = in_1[247] + e1[0][247] %3329;
                                                                                                                                                                                 u[0][248] = in_1[248] + e1[0][248] %3329;
                                                                                                                                                                                 u[0][249] = in_1[249] + e1[0][249] %3329;
                                                                                                                                                                                 u[0][250] = in_1[250] + e1[0][250] %3329;
                                                                                                                                                                                 u[0][251] = in_1[251] + e1[0][251] %3329;
                                                                                                                                                                                 u[0][252] = in_1[252] + e1[0][252] %3329;
                                                                                                                                                                                 u[0][253] = in_1[253] + e1[0][253] %3329;
                                                                                                                                                                                 u[0][254] = in_1[254] + e1[0][254] %3329;
                                                                                                                                                                                 u[0][255] = in_1[255] + e1[0][255] %3329;
                                                                                                                                                                                 u[1][0] = in_2[0] + e1[1][0] %3329;
                                                                                                                                                                                 u[1][1] = in_2[1] + e1[1][1] %3329;
                                                                                                                                                                                 u[1][2] = in_2[2] + e1[1][2] %3329;
                                                                                                                                                                                 u[1][3] = in_2[3] + e1[1][3] %3329;
                                                                                                                                                                                 u[1][4] = in_2[4] + e1[1][4] %3329;
                                                                                                                                                                                 u[1][5] = in_2[5] + e1[1][5] %3329;
                                                                                                                                                                                 u[1][6] = in_2[6] + e1[1][6] %3329;
                                                                                                                                                                                 u[1][7] = in_2[7] + e1[1][7] %3329;
                                                                                                                                                                                 u[1][8] = in_2[8] + e1[1][8] %3329;
                                                                                                                                                                                 u[1][9] = in_2[9] + e1[1][9] %3329;
                                                                                                                                                                                 u[1][10] = in_2[10] + e1[1][10] %3329;
                                                                                                                                                                                 u[1][11] = in_2[11] + e1[1][11] %3329;
                                                                                                                                                                                 u[1][12] = in_2[12] + e1[1][12] %3329;
                                                                                                                                                                                 u[1][13] = in_2[13] + e1[1][13] %3329;
                                                                                                                                                                                 u[1][14] = in_2[14] + e1[1][14] %3329;
                                                                                                                                                                                 u[1][15] = in_2[15] + e1[1][15] %3329;
                                                                                                                                                                                 u[1][16] = in_2[16] + e1[1][16] %3329;
                                                                                                                                                                                 u[1][17] = in_2[17] + e1[1][17] %3329;
                                                                                                                                                                                 u[1][18] = in_2[18] + e1[1][18] %3329;
                                                                                                                                                                                 u[1][19] = in_2[19] + e1[1][19] %3329;
                                                                                                                                                                                 u[1][20] = in_2[20] + e1[1][20] %3329;
                                                                                                                                                                                 u[1][21] = in_2[21] + e1[1][21] %3329;
                                                                                                                                                                                 u[1][22] = in_2[22] + e1[1][22] %3329;
                                                                                                                                                                                 u[1][23] = in_2[23] + e1[1][23] %3329;
                                                                                                                                                                                 u[1][24] = in_2[24] + e1[1][24] %3329;
                                                                                                                                                                                 u[1][25] = in_2[25] + e1[1][25] %3329;
                                                                                                                                                                                 u[1][26] = in_2[26] + e1[1][26] %3329;
                                                                                                                                                                                 u[1][27] = in_2[27] + e1[1][27] %3329;
                                                                                                                                                                                 u[1][28] = in_2[28] + e1[1][28] %3329;
                                                                                                                                                                                 u[1][29] = in_2[29] + e1[1][29] %3329;
                                                                                                                                                                                 u[1][30] = in_2[30] + e1[1][30] %3329;
                                                                                                                                                                                 u[1][31] = in_2[31] + e1[1][31] %3329;
                                                                                                                                                                                 u[1][32] = in_2[32] + e1[1][32] %3329;
                                                                                                                                                                                 u[1][33] = in_2[33] + e1[1][33] %3329;
                                                                                                                                                                                 u[1][34] = in_2[34] + e1[1][34] %3329;
                                                                                                                                                                                 u[1][35] = in_2[35] + e1[1][35] %3329;
                                                                                                                                                                                 u[1][36] = in_2[36] + e1[1][36] %3329;
                                                                                                                                                                                 u[1][37] = in_2[37] + e1[1][37] %3329;
                                                                                                                                                                                 u[1][38] = in_2[38] + e1[1][38] %3329;
                                                                                                                                                                                 u[1][39] = in_2[39] + e1[1][39] %3329;
                                                                                                                                                                                 u[1][40] = in_2[40] + e1[1][40] %3329;
                                                                                                                                                                                 u[1][41] = in_2[41] + e1[1][41] %3329;
                                                                                                                                                                                 u[1][42] = in_2[42] + e1[1][42] %3329;
                                                                                                                                                                                 u[1][43] = in_2[43] + e1[1][43] %3329;
                                                                                                                                                                                 u[1][44] = in_2[44] + e1[1][44] %3329;
                                                                                                                                                                                 u[1][45] = in_2[45] + e1[1][45] %3329;
                                                                                                                                                                                 u[1][46] = in_2[46] + e1[1][46] %3329;
                                                                                                                                                                                 u[1][47] = in_2[47] + e1[1][47] %3329;
                                                                                                                                                                                 u[1][48] = in_2[48] + e1[1][48] %3329;
                                                                                                                                                                                 u[1][49] = in_2[49] + e1[1][49] %3329;
                                                                                                                                                                                 u[1][50] = in_2[50] + e1[1][50] %3329;
                                                                                                                                                                                 u[1][51] = in_2[51] + e1[1][51] %3329;
                                                                                                                                                                                 u[1][52] = in_2[52] + e1[1][52] %3329;
                                                                                                                                                                                 u[1][53] = in_2[53] + e1[1][53] %3329;
                                                                                                                                                                                 u[1][54] = in_2[54] + e1[1][54] %3329;
                                                                                                                                                                                 u[1][55] = in_2[55] + e1[1][55] %3329;
                                                                                                                                                                                 u[1][56] = in_2[56] + e1[1][56] %3329;
                                                                                                                                                                                 u[1][57] = in_2[57] + e1[1][57] %3329;
                                                                                                                                                                                 u[1][58] = in_2[58] + e1[1][58] %3329;
                                                                                                                                                                                 u[1][59] = in_2[59] + e1[1][59] %3329;
                                                                                                                                                                                 u[1][60] = in_2[60] + e1[1][60] %3329;
                                                                                                                                                                                 u[1][61] = in_2[61] + e1[1][61] %3329;
                                                                                                                                                                                 u[1][62] = in_2[62] + e1[1][62] %3329;
                                                                                                                                                                                 u[1][63] = in_2[63] + e1[1][63] %3329;
                                                                                                                                                                                 u[1][64] = in_2[64] + e1[1][64] %3329;
                                                                                                                                                                                 u[1][65] = in_2[65] + e1[1][65] %3329;
                                                                                                                                                                                 u[1][66] = in_2[66] + e1[1][66] %3329;
                                                                                                                                                                                 u[1][67] = in_2[67] + e1[1][67] %3329;
                                                                                                                                                                                 u[1][68] = in_2[68] + e1[1][68] %3329;
                                                                                                                                                                                 u[1][69] = in_2[69] + e1[1][69] %3329;
                                                                                                                                                                                 u[1][70] = in_2[70] + e1[1][70] %3329;
                                                                                                                                                                                 u[1][71] = in_2[71] + e1[1][71] %3329;
                                                                                                                                                                                 u[1][72] = in_2[72] + e1[1][72] %3329;
                                                                                                                                                                                 u[1][73] = in_2[73] + e1[1][73] %3329;
                                                                                                                                                                                 u[1][74] = in_2[74] + e1[1][74] %3329;
                                                                                                                                                                                 u[1][75] = in_2[75] + e1[1][75] %3329;
                                                                                                                                                                                 u[1][76] = in_2[76] + e1[1][76] %3329;
                                                                                                                                                                                 u[1][77] = in_2[77] + e1[1][77] %3329;
                                                                                                                                                                                 u[1][78] = in_2[78] + e1[1][78] %3329;
                                                                                                                                                                                 u[1][79] = in_2[79] + e1[1][79] %3329;
                                                                                                                                                                                 u[1][80] = in_2[80] + e1[1][80] %3329;
                                                                                                                                                                                 u[1][81] = in_2[81] + e1[1][81] %3329;
                                                                                                                                                                                 u[1][82] = in_2[82] + e1[1][82] %3329;
                                                                                                                                                                                 u[1][83] = in_2[83] + e1[1][83] %3329;
                                                                                                                                                                                 u[1][84] = in_2[84] + e1[1][84] %3329;
                                                                                                                                                                                 u[1][85] = in_2[85] + e1[1][85] %3329;
                                                                                                                                                                                 u[1][86] = in_2[86] + e1[1][86] %3329;
                                                                                                                                                                                 u[1][87] = in_2[87] + e1[1][87] %3329;
                                                                                                                                                                                 u[1][88] = in_2[88] + e1[1][88] %3329;
                                                                                                                                                                                 u[1][89] = in_2[89] + e1[1][89] %3329;
                                                                                                                                                                                 u[1][90] = in_2[90] + e1[1][90] %3329;
                                                                                                                                                                                 u[1][91] = in_2[91] + e1[1][91] %3329;
                                                                                                                                                                                 u[1][92] = in_2[92] + e1[1][92] %3329;
                                                                                                                                                                                 u[1][93] = in_2[93] + e1[1][93] %3329;
                                                                                                                                                                                 u[1][94] = in_2[94] + e1[1][94] %3329;
                                                                                                                                                                                 u[1][95] = in_2[95] + e1[1][95] %3329;
                                                                                                                                                                                 u[1][96] = in_2[96] + e1[1][96] %3329;
                                                                                                                                                                                 u[1][97] = in_2[97] + e1[1][97] %3329;
                                                                                                                                                                                 u[1][98] = in_2[98] + e1[1][98] %3329;
                                                                                                                                                                                 u[1][99] = in_2[99] + e1[1][99] %3329;
                                                                                                                                                                                 u[1][100] = in_2[100] + e1[1][100] %3329;
                                                                                                                                                                                 u[1][101] = in_2[101] + e1[1][101] %3329;
                                                                                                                                                                                 u[1][102] = in_2[102] + e1[1][102] %3329;
                                                                                                                                                                                 u[1][103] = in_2[103] + e1[1][103] %3329;
                                                                                                                                                                                 u[1][104] = in_2[104] + e1[1][104] %3329;
                                                                                                                                                                                 u[1][105] = in_2[105] + e1[1][105] %3329;
                                                                                                                                                                                 u[1][106] = in_2[106] + e1[1][106] %3329;
                                                                                                                                                                                 u[1][107] = in_2[107] + e1[1][107] %3329;
                                                                                                                                                                                 u[1][108] = in_2[108] + e1[1][108] %3329;
                                                                                                                                                                                 u[1][109] = in_2[109] + e1[1][109] %3329;
                                                                                                                                                                                 u[1][110] = in_2[110] + e1[1][110] %3329;
                                                                                                                                                                                 u[1][111] = in_2[111] + e1[1][111] %3329;
                                                                                                                                                                                 u[1][112] = in_2[112] + e1[1][112] %3329;
                                                                                                                                                                                 u[1][113] = in_2[113] + e1[1][113] %3329;
                                                                                                                                                                                 u[1][114] = in_2[114] + e1[1][114] %3329;
                                                                                                                                                                                 u[1][115] = in_2[115] + e1[1][115] %3329;
                                                                                                                                                                                 u[1][116] = in_2[116] + e1[1][116] %3329;
                                                                                                                                                                                 u[1][117] = in_2[117] + e1[1][117] %3329;
                                                                                                                                                                                 u[1][118] = in_2[118] + e1[1][118] %3329;
                                                                                                                                                                                 u[1][119] = in_2[119] + e1[1][119] %3329;
                                                                                                                                                                                 u[1][120] = in_2[120] + e1[1][120] %3329;
                                                                                                                                                                                 u[1][121] = in_2[121] + e1[1][121] %3329;
                                                                                                                                                                                 u[1][122] = in_2[122] + e1[1][122] %3329;
                                                                                                                                                                                 u[1][123] = in_2[123] + e1[1][123] %3329;
                                                                                                                                                                                 u[1][124] = in_2[124] + e1[1][124] %3329;
                                                                                                                                                                                 u[1][125] = in_2[125] + e1[1][125] %3329;
                                                                                                                                                                                 u[1][126] = in_2[126] + e1[1][126] %3329;
                                                                                                                                                                                 u[1][127] = in_2[127] + e1[1][127] %3329;
                                                                                                                                                                                 u[1][128] = in_2[128] + e1[1][128] %3329;
                                                                                                                                                                                 u[1][129] = in_2[129] + e1[1][129] %3329;
                                                                                                                                                                                 u[1][130] = in_2[130] + e1[1][130] %3329;
                                                                                                                                                                                 u[1][131] = in_2[131] + e1[1][131] %3329;
                                                                                                                                                                                 u[1][132] = in_2[132] + e1[1][132] %3329;
                                                                                                                                                                                 u[1][133] = in_2[133] + e1[1][133] %3329;
                                                                                                                                                                                 u[1][134] = in_2[134] + e1[1][134] %3329;
                                                                                                                                                                                 u[1][135] = in_2[135] + e1[1][135] %3329;
                                                                                                                                                                                 u[1][136] = in_2[136] + e1[1][136] %3329;
                                                                                                                                                                                 u[1][137] = in_2[137] + e1[1][137] %3329;
                                                                                                                                                                                 u[1][138] = in_2[138] + e1[1][138] %3329;
                                                                                                                                                                                 u[1][139] = in_2[139] + e1[1][139] %3329;
                                                                                                                                                                                 u[1][140] = in_2[140] + e1[1][140] %3329;
                                                                                                                                                                                 u[1][141] = in_2[141] + e1[1][141] %3329;
                                                                                                                                                                                 u[1][142] = in_2[142] + e1[1][142] %3329;
                                                                                                                                                                                 u[1][143] = in_2[143] + e1[1][143] %3329;
                                                                                                                                                                                 u[1][144] = in_2[144] + e1[1][144] %3329;
                                                                                                                                                                                 u[1][145] = in_2[145] + e1[1][145] %3329;
                                                                                                                                                                                 u[1][146] = in_2[146] + e1[1][146] %3329;
                                                                                                                                                                                 u[1][147] = in_2[147] + e1[1][147] %3329;
                                                                                                                                                                                 u[1][148] = in_2[148] + e1[1][148] %3329;
                                                                                                                                                                                 u[1][149] = in_2[149] + e1[1][149] %3329;
                                                                                                                                                                                 u[1][150] = in_2[150] + e1[1][150] %3329;
                                                                                                                                                                                 u[1][151] = in_2[151] + e1[1][151] %3329;
                                                                                                                                                                                 u[1][152] = in_2[152] + e1[1][152] %3329;
                                                                                                                                                                                 u[1][153] = in_2[153] + e1[1][153] %3329;
                                                                                                                                                                                 u[1][154] = in_2[154] + e1[1][154] %3329;
                                                                                                                                                                                 u[1][155] = in_2[155] + e1[1][155] %3329;
                                                                                                                                                                                 u[1][156] = in_2[156] + e1[1][156] %3329;
                                                                                                                                                                                 u[1][157] = in_2[157] + e1[1][157] %3329;
                                                                                                                                                                                 u[1][158] = in_2[158] + e1[1][158] %3329;
                                                                                                                                                                                 u[1][159] = in_2[159] + e1[1][159] %3329;
                                                                                                                                                                                 u[1][160] = in_2[160] + e1[1][160] %3329;
                                                                                                                                                                                 u[1][161] = in_2[161] + e1[1][161] %3329;
                                                                                                                                                                                 u[1][162] = in_2[162] + e1[1][162] %3329;
                                                                                                                                                                                 u[1][163] = in_2[163] + e1[1][163] %3329;
                                                                                                                                                                                 u[1][164] = in_2[164] + e1[1][164] %3329;
                                                                                                                                                                                 u[1][165] = in_2[165] + e1[1][165] %3329;
                                                                                                                                                                                 u[1][166] = in_2[166] + e1[1][166] %3329;
                                                                                                                                                                                 u[1][167] = in_2[167] + e1[1][167] %3329;
                                                                                                                                                                                 u[1][168] = in_2[168] + e1[1][168] %3329;
                                                                                                                                                                                 u[1][169] = in_2[169] + e1[1][169] %3329;
                                                                                                                                                                                 u[1][170] = in_2[170] + e1[1][170] %3329;
                                                                                                                                                                                 u[1][171] = in_2[171] + e1[1][171] %3329;
                                                                                                                                                                                 u[1][172] = in_2[172] + e1[1][172] %3329;
                                                                                                                                                                                 u[1][173] = in_2[173] + e1[1][173] %3329;
                                                                                                                                                                                 u[1][174] = in_2[174] + e1[1][174] %3329;
                                                                                                                                                                                 u[1][175] = in_2[175] + e1[1][175] %3329;
                                                                                                                                                                                 u[1][176] = in_2[176] + e1[1][176] %3329;
                                                                                                                                                                                 u[1][177] = in_2[177] + e1[1][177] %3329;
                                                                                                                                                                                 u[1][178] = in_2[178] + e1[1][178] %3329;
                                                                                                                                                                                 u[1][179] = in_2[179] + e1[1][179] %3329;
                                                                                                                                                                                 u[1][180] = in_2[180] + e1[1][180] %3329;
                                                                                                                                                                                 u[1][181] = in_2[181] + e1[1][181] %3329;
                                                                                                                                                                                 u[1][182] = in_2[182] + e1[1][182] %3329;
                                                                                                                                                                                 u[1][183] = in_2[183] + e1[1][183] %3329;
                                                                                                                                                                                 u[1][184] = in_2[184] + e1[1][184] %3329;
                                                                                                                                                                                 u[1][185] = in_2[185] + e1[1][185] %3329;
                                                                                                                                                                                 u[1][186] = in_2[186] + e1[1][186] %3329;
                                                                                                                                                                                 u[1][187] = in_2[187] + e1[1][187] %3329;
                                                                                                                                                                                 u[1][188] = in_2[188] + e1[1][188] %3329;
                                                                                                                                                                                 u[1][189] = in_2[189] + e1[1][189] %3329;
                                                                                                                                                                                 u[1][190] = in_2[190] + e1[1][190] %3329;
                                                                                                                                                                                 u[1][191] = in_2[191] + e1[1][191] %3329;
                                                                                                                                                                                 u[1][192] = in_2[192] + e1[1][192] %3329;
                                                                                                                                                                                 u[1][193] = in_2[193] + e1[1][193] %3329;
                                                                                                                                                                                 u[1][194] = in_2[194] + e1[1][194] %3329;
                                                                                                                                                                                 u[1][195] = in_2[195] + e1[1][195] %3329;
                                                                                                                                                                                 u[1][196] = in_2[196] + e1[1][196] %3329;
                                                                                                                                                                                 u[1][197] = in_2[197] + e1[1][197] %3329;
                                                                                                                                                                                 u[1][198] = in_2[198] + e1[1][198] %3329;
                                                                                                                                                                                 u[1][199] = in_2[199] + e1[1][199] %3329;
                                                                                                                                                                                 u[1][200] = in_2[200] + e1[1][200] %3329;
                                                                                                                                                                                 u[1][201] = in_2[201] + e1[1][201] %3329;
                                                                                                                                                                                 u[1][202] = in_2[202] + e1[1][202] %3329;
                                                                                                                                                                                 u[1][203] = in_2[203] + e1[1][203] %3329;
                                                                                                                                                                                 u[1][204] = in_2[204] + e1[1][204] %3329;
                                                                                                                                                                                 u[1][205] = in_2[205] + e1[1][205] %3329;
                                                                                                                                                                                 u[1][206] = in_2[206] + e1[1][206] %3329;
                                                                                                                                                                                 u[1][207] = in_2[207] + e1[1][207] %3329;
                                                                                                                                                                                 u[1][208] = in_2[208] + e1[1][208] %3329;
                                                                                                                                                                                 u[1][209] = in_2[209] + e1[1][209] %3329;
                                                                                                                                                                                 u[1][210] = in_2[210] + e1[1][210] %3329;
                                                                                                                                                                                 u[1][211] = in_2[211] + e1[1][211] %3329;
                                                                                                                                                                                 u[1][212] = in_2[212] + e1[1][212] %3329;
                                                                                                                                                                                 u[1][213] = in_2[213] + e1[1][213] %3329;
                                                                                                                                                                                 u[1][214] = in_2[214] + e1[1][214] %3329;
                                                                                                                                                                                 u[1][215] = in_2[215] + e1[1][215] %3329;
                                                                                                                                                                                 u[1][216] = in_2[216] + e1[1][216] %3329;
                                                                                                                                                                                 u[1][217] = in_2[217] + e1[1][217] %3329;
                                                                                                                                                                                 u[1][218] = in_2[218] + e1[1][218] %3329;
                                                                                                                                                                                 u[1][219] = in_2[219] + e1[1][219] %3329;
                                                                                                                                                                                 u[1][220] = in_2[220] + e1[1][220] %3329;
                                                                                                                                                                                 u[1][221] = in_2[221] + e1[1][221] %3329;
                                                                                                                                                                                 u[1][222] = in_2[222] + e1[1][222] %3329;
                                                                                                                                                                                 u[1][223] = in_2[223] + e1[1][223] %3329;
                                                                                                                                                                                 u[1][224] = in_2[224] + e1[1][224] %3329;
                                                                                                                                                                                 u[1][225] = in_2[225] + e1[1][225] %3329;
                                                                                                                                                                                 u[1][226] = in_2[226] + e1[1][226] %3329;
                                                                                                                                                                                 u[1][227] = in_2[227] + e1[1][227] %3329;
                                                                                                                                                                                 u[1][228] = in_2[228] + e1[1][228] %3329;
                                                                                                                                                                                 u[1][229] = in_2[229] + e1[1][229] %3329;
                                                                                                                                                                                 u[1][230] = in_2[230] + e1[1][230] %3329;
                                                                                                                                                                                 u[1][231] = in_2[231] + e1[1][231] %3329;
                                                                                                                                                                                 u[1][232] = in_2[232] + e1[1][232] %3329;
                                                                                                                                                                                 u[1][233] = in_2[233] + e1[1][233] %3329;
                                                                                                                                                                                 u[1][234] = in_2[234] + e1[1][234] %3329;
                                                                                                                                                                                 u[1][235] = in_2[235] + e1[1][235] %3329;
                                                                                                                                                                                 u[1][236] = in_2[236] + e1[1][236] %3329;
                                                                                                                                                                                 u[1][237] = in_2[237] + e1[1][237] %3329;
                                                                                                                                                                                 u[1][238] = in_2[238] + e1[1][238] %3329;
                                                                                                                                                                                 u[1][239] = in_2[239] + e1[1][239] %3329;
                                                                                                                                                                                 u[1][240] = in_2[240] + e1[1][240] %3329;
                                                                                                                                                                                 u[1][241] = in_2[241] + e1[1][241] %3329;
                                                                                                                                                                                 u[1][242] = in_2[242] + e1[1][242] %3329;
                                                                                                                                                                                 u[1][243] = in_2[243] + e1[1][243] %3329;
                                                                                                                                                                                 u[1][244] = in_2[244] + e1[1][244] %3329;
                                                                                                                                                                                 u[1][245] = in_2[245] + e1[1][245] %3329;
                                                                                                                                                                                 u[1][246] = in_2[246] + e1[1][246] %3329;
                                                                                                                                                                                 u[1][247] = in_2[247] + e1[1][247] %3329;
                                                                                                                                                                                 u[1][248] = in_2[248] + e1[1][248] %3329;
                                                                                                                                                                                 u[1][249] = in_2[249] + e1[1][249] %3329;
                                                                                                                                                                                 u[1][250] = in_2[250] + e1[1][250] %3329;
                                                                                                                                                                                 u[1][251] = in_2[251] + e1[1][251] %3329;
                                                                                                                                                                                 u[1][252] = in_2[252] + e1[1][252] %3329;
                                                                                                                                                                                 u[1][253] = in_2[253] + e1[1][253] %3329;
                                                                                                                                                                                 u[1][254] = in_2[254] + e1[1][254] %3329;
                                                                                                                                                                                 u[1][255] = in_2[255] + e1[1][255] %3329;
                                                                                                                                                                                 u[2][0] = in_3[0] + e1[2][0] %3329;
                                                                                                                                                                                 u[2][1] = in_3[1] + e1[2][1] %3329;
                                                                                                                                                                                 u[2][2] = in_3[2] + e1[2][2] %3329;
                                                                                                                                                                                 u[2][3] = in_3[3] + e1[2][3] %3329;
                                                                                                                                                                                 u[2][4] = in_3[4] + e1[2][4] %3329;
                                                                                                                                                                                 u[2][5] = in_3[5] + e1[2][5] %3329;
                                                                                                                                                                                 u[2][6] = in_3[6] + e1[2][6] %3329;
                                                                                                                                                                                 u[2][7] = in_3[7] + e1[2][7] %3329;
                                                                                                                                                                                 u[2][8] = in_3[8] + e1[2][8] %3329;
                                                                                                                                                                                 u[2][9] = in_3[9] + e1[2][9] %3329;
                                                                                                                                                                                 u[2][10] = in_3[10] + e1[2][10] %3329;
                                                                                                                                                                                 u[2][11] = in_3[11] + e1[2][11] %3329;
                                                                                                                                                                                 u[2][12] = in_3[12] + e1[2][12] %3329;
                                                                                                                                                                                 u[2][13] = in_3[13] + e1[2][13] %3329;
                                                                                                                                                                                 u[2][14] = in_3[14] + e1[2][14] %3329;
                                                                                                                                                                                 u[2][15] = in_3[15] + e1[2][15] %3329;
                                                                                                                                                                                 u[2][16] = in_3[16] + e1[2][16] %3329;
                                                                                                                                                                                 u[2][17] = in_3[17] + e1[2][17] %3329;
                                                                                                                                                                                 u[2][18] = in_3[18] + e1[2][18] %3329;
                                                                                                                                                                                 u[2][19] = in_3[19] + e1[2][19] %3329;
                                                                                                                                                                                 u[2][20] = in_3[20] + e1[2][20] %3329;
                                                                                                                                                                                 u[2][21] = in_3[21] + e1[2][21] %3329;
                                                                                                                                                                                 u[2][22] = in_3[22] + e1[2][22] %3329;
                                                                                                                                                                                 u[2][23] = in_3[23] + e1[2][23] %3329;
                                                                                                                                                                                 u[2][24] = in_3[24] + e1[2][24] %3329;
                                                                                                                                                                                 u[2][25] = in_3[25] + e1[2][25] %3329;
                                                                                                                                                                                 u[2][26] = in_3[26] + e1[2][26] %3329;
                                                                                                                                                                                 u[2][27] = in_3[27] + e1[2][27] %3329;
                                                                                                                                                                                 u[2][28] = in_3[28] + e1[2][28] %3329;
                                                                                                                                                                                 u[2][29] = in_3[29] + e1[2][29] %3329;
                                                                                                                                                                                 u[2][30] = in_3[30] + e1[2][30] %3329;
                                                                                                                                                                                 u[2][31] = in_3[31] + e1[2][31] %3329;
                                                                                                                                                                                 u[2][32] = in_3[32] + e1[2][32] %3329;
                                                                                                                                                                                 u[2][33] = in_3[33] + e1[2][33] %3329;
                                                                                                                                                                                 u[2][34] = in_3[34] + e1[2][34] %3329;
                                                                                                                                                                                 u[2][35] = in_3[35] + e1[2][35] %3329;
                                                                                                                                                                                 u[2][36] = in_3[36] + e1[2][36] %3329;
                                                                                                                                                                                 u[2][37] = in_3[37] + e1[2][37] %3329;
                                                                                                                                                                                 u[2][38] = in_3[38] + e1[2][38] %3329;
                                                                                                                                                                                 u[2][39] = in_3[39] + e1[2][39] %3329;
                                                                                                                                                                                 u[2][40] = in_3[40] + e1[2][40] %3329;
                                                                                                                                                                                 u[2][41] = in_3[41] + e1[2][41] %3329;
                                                                                                                                                                                 u[2][42] = in_3[42] + e1[2][42] %3329;
                                                                                                                                                                                 u[2][43] = in_3[43] + e1[2][43] %3329;
                                                                                                                                                                                 u[2][44] = in_3[44] + e1[2][44] %3329;
                                                                                                                                                                                 u[2][45] = in_3[45] + e1[2][45] %3329;
                                                                                                                                                                                 u[2][46] = in_3[46] + e1[2][46] %3329;
                                                                                                                                                                                 u[2][47] = in_3[47] + e1[2][47] %3329;
                                                                                                                                                                                 u[2][48] = in_3[48] + e1[2][48] %3329;
                                                                                                                                                                                 u[2][49] = in_3[49] + e1[2][49] %3329;
                                                                                                                                                                                 u[2][50] = in_3[50] + e1[2][50] %3329;
                                                                                                                                                                                 u[2][51] = in_3[51] + e1[2][51] %3329;
                                                                                                                                                                                 u[2][52] = in_3[52] + e1[2][52] %3329;
                                                                                                                                                                                 u[2][53] = in_3[53] + e1[2][53] %3329;
                                                                                                                                                                                 u[2][54] = in_3[54] + e1[2][54] %3329;
                                                                                                                                                                                 u[2][55] = in_3[55] + e1[2][55] %3329;
                                                                                                                                                                                 u[2][56] = in_3[56] + e1[2][56] %3329;
                                                                                                                                                                                 u[2][57] = in_3[57] + e1[2][57] %3329;
                                                                                                                                                                                 u[2][58] = in_3[58] + e1[2][58] %3329;
                                                                                                                                                                                 u[2][59] = in_3[59] + e1[2][59] %3329;
                                                                                                                                                                                 u[2][60] = in_3[60] + e1[2][60] %3329;
                                                                                                                                                                                 u[2][61] = in_3[61] + e1[2][61] %3329;
                                                                                                                                                                                 u[2][62] = in_3[62] + e1[2][62] %3329;
                                                                                                                                                                                 u[2][63] = in_3[63] + e1[2][63] %3329;
                                                                                                                                                                                 u[2][64] = in_3[64] + e1[2][64] %3329;
                                                                                                                                                                                 u[2][65] = in_3[65] + e1[2][65] %3329;
                                                                                                                                                                                 u[2][66] = in_3[66] + e1[2][66] %3329;
                                                                                                                                                                                 u[2][67] = in_3[67] + e1[2][67] %3329;
                                                                                                                                                                                 u[2][68] = in_3[68] + e1[2][68] %3329;
                                                                                                                                                                                 u[2][69] = in_3[69] + e1[2][69] %3329;
                                                                                                                                                                                 u[2][70] = in_3[70] + e1[2][70] %3329;
                                                                                                                                                                                 u[2][71] = in_3[71] + e1[2][71] %3329;
                                                                                                                                                                                 u[2][72] = in_3[72] + e1[2][72] %3329;
                                                                                                                                                                                 u[2][73] = in_3[73] + e1[2][73] %3329;
                                                                                                                                                                                 u[2][74] = in_3[74] + e1[2][74] %3329;
                                                                                                                                                                                 u[2][75] = in_3[75] + e1[2][75] %3329;
                                                                                                                                                                                 u[2][76] = in_3[76] + e1[2][76] %3329;
                                                                                                                                                                                 u[2][77] = in_3[77] + e1[2][77] %3329;
                                                                                                                                                                                 u[2][78] = in_3[78] + e1[2][78] %3329;
                                                                                                                                                                                 u[2][79] = in_3[79] + e1[2][79] %3329;
                                                                                                                                                                                 u[2][80] = in_3[80] + e1[2][80] %3329;
                                                                                                                                                                                 u[2][81] = in_3[81] + e1[2][81] %3329;
                                                                                                                                                                                 u[2][82] = in_3[82] + e1[2][82] %3329;
                                                                                                                                                                                 u[2][83] = in_3[83] + e1[2][83] %3329;
                                                                                                                                                                                 u[2][84] = in_3[84] + e1[2][84] %3329;
                                                                                                                                                                                 u[2][85] = in_3[85] + e1[2][85] %3329;
                                                                                                                                                                                 u[2][86] = in_3[86] + e1[2][86] %3329;
                                                                                                                                                                                 u[2][87] = in_3[87] + e1[2][87] %3329;
                                                                                                                                                                                 u[2][88] = in_3[88] + e1[2][88] %3329;
                                                                                                                                                                                 u[2][89] = in_3[89] + e1[2][89] %3329;
                                                                                                                                                                                 u[2][90] = in_3[90] + e1[2][90] %3329;
                                                                                                                                                                                 u[2][91] = in_3[91] + e1[2][91] %3329;
                                                                                                                                                                                 u[2][92] = in_3[92] + e1[2][92] %3329;
                                                                                                                                                                                 u[2][93] = in_3[93] + e1[2][93] %3329;
                                                                                                                                                                                 u[2][94] = in_3[94] + e1[2][94] %3329;
                                                                                                                                                                                 u[2][95] = in_3[95] + e1[2][95] %3329;
                                                                                                                                                                                 u[2][96] = in_3[96] + e1[2][96] %3329;
                                                                                                                                                                                 u[2][97] = in_3[97] + e1[2][97] %3329;
                                                                                                                                                                                 u[2][98] = in_3[98] + e1[2][98] %3329;
                                                                                                                                                                                 u[2][99] = in_3[99] + e1[2][99] %3329;
                                                                                                                                                                                 u[2][100] = in_3[100] + e1[2][100] %3329;
                                                                                                                                                                                 u[2][101] = in_3[101] + e1[2][101] %3329;
                                                                                                                                                                                 u[2][102] = in_3[102] + e1[2][102] %3329;
                                                                                                                                                                                 u[2][103] = in_3[103] + e1[2][103] %3329;
                                                                                                                                                                                 u[2][104] = in_3[104] + e1[2][104] %3329;
                                                                                                                                                                                 u[2][105] = in_3[105] + e1[2][105] %3329;
                                                                                                                                                                                 u[2][106] = in_3[106] + e1[2][106] %3329;
                                                                                                                                                                                 u[2][107] = in_3[107] + e1[2][107] %3329;
                                                                                                                                                                                 u[2][108] = in_3[108] + e1[2][108] %3329;
                                                                                                                                                                                 u[2][109] = in_3[109] + e1[2][109] %3329;
                                                                                                                                                                                 u[2][110] = in_3[110] + e1[2][110] %3329;
                                                                                                                                                                                 u[2][111] = in_3[111] + e1[2][111] %3329;
                                                                                                                                                                                 u[2][112] = in_3[112] + e1[2][112] %3329;
                                                                                                                                                                                 u[2][113] = in_3[113] + e1[2][113] %3329;
                                                                                                                                                                                 u[2][114] = in_3[114] + e1[2][114] %3329;
                                                                                                                                                                                 u[2][115] = in_3[115] + e1[2][115] %3329;
                                                                                                                                                                                 u[2][116] = in_3[116] + e1[2][116] %3329;
                                                                                                                                                                                 u[2][117] = in_3[117] + e1[2][117] %3329;
                                                                                                                                                                                 u[2][118] = in_3[118] + e1[2][118] %3329;
                                                                                                                                                                                 u[2][119] = in_3[119] + e1[2][119] %3329;
                                                                                                                                                                                 u[2][120] = in_3[120] + e1[2][120] %3329;
                                                                                                                                                                                 u[2][121] = in_3[121] + e1[2][121] %3329;
                                                                                                                                                                                 u[2][122] = in_3[122] + e1[2][122] %3329;
                                                                                                                                                                                 u[2][123] = in_3[123] + e1[2][123] %3329;
                                                                                                                                                                                 u[2][124] = in_3[124] + e1[2][124] %3329;
                                                                                                                                                                                 u[2][125] = in_3[125] + e1[2][125] %3329;
                                                                                                                                                                                 u[2][126] = in_3[126] + e1[2][126] %3329;
                                                                                                                                                                                 u[2][127] = in_3[127] + e1[2][127] %3329;
                                                                                                                                                                                 u[2][128] = in_3[128] + e1[2][128] %3329;
                                                                                                                                                                                 u[2][129] = in_3[129] + e1[2][129] %3329;
                                                                                                                                                                                 u[2][130] = in_3[130] + e1[2][130] %3329;
                                                                                                                                                                                 u[2][131] = in_3[131] + e1[2][131] %3329;
                                                                                                                                                                                 u[2][132] = in_3[132] + e1[2][132] %3329;
                                                                                                                                                                                 u[2][133] = in_3[133] + e1[2][133] %3329;
                                                                                                                                                                                 u[2][134] = in_3[134] + e1[2][134] %3329;
                                                                                                                                                                                 u[2][135] = in_3[135] + e1[2][135] %3329;
                                                                                                                                                                                 u[2][136] = in_3[136] + e1[2][136] %3329;
                                                                                                                                                                                 u[2][137] = in_3[137] + e1[2][137] %3329;
                                                                                                                                                                                 u[2][138] = in_3[138] + e1[2][138] %3329;
                                                                                                                                                                                 u[2][139] = in_3[139] + e1[2][139] %3329;
                                                                                                                                                                                 u[2][140] = in_3[140] + e1[2][140] %3329;
                                                                                                                                                                                 u[2][141] = in_3[141] + e1[2][141] %3329;
                                                                                                                                                                                 u[2][142] = in_3[142] + e1[2][142] %3329;
                                                                                                                                                                                 u[2][143] = in_3[143] + e1[2][143] %3329;
                                                                                                                                                                                 u[2][144] = in_3[144] + e1[2][144] %3329;
                                                                                                                                                                                 u[2][145] = in_3[145] + e1[2][145] %3329;
                                                                                                                                                                                 u[2][146] = in_3[146] + e1[2][146] %3329;
                                                                                                                                                                                 u[2][147] = in_3[147] + e1[2][147] %3329;
                                                                                                                                                                                 u[2][148] = in_3[148] + e1[2][148] %3329;
                                                                                                                                                                                 u[2][149] = in_3[149] + e1[2][149] %3329;
                                                                                                                                                                                 u[2][150] = in_3[150] + e1[2][150] %3329;
                                                                                                                                                                                 u[2][151] = in_3[151] + e1[2][151] %3329;
                                                                                                                                                                                 u[2][152] = in_3[152] + e1[2][152] %3329;
                                                                                                                                                                                 u[2][153] = in_3[153] + e1[2][153] %3329;
                                                                                                                                                                                 u[2][154] = in_3[154] + e1[2][154] %3329;
                                                                                                                                                                                 u[2][155] = in_3[155] + e1[2][155] %3329;
                                                                                                                                                                                 u[2][156] = in_3[156] + e1[2][156] %3329;
                                                                                                                                                                                 u[2][157] = in_3[157] + e1[2][157] %3329;
                                                                                                                                                                                 u[2][158] = in_3[158] + e1[2][158] %3329;
                                                                                                                                                                                 u[2][159] = in_3[159] + e1[2][159] %3329;
                                                                                                                                                                                 u[2][160] = in_3[160] + e1[2][160] %3329;
                                                                                                                                                                                 u[2][161] = in_3[161] + e1[2][161] %3329;
                                                                                                                                                                                 u[2][162] = in_3[162] + e1[2][162] %3329;
                                                                                                                                                                                 u[2][163] = in_3[163] + e1[2][163] %3329;
                                                                                                                                                                                 u[2][164] = in_3[164] + e1[2][164] %3329;
                                                                                                                                                                                 u[2][165] = in_3[165] + e1[2][165] %3329;
                                                                                                                                                                                 u[2][166] = in_3[166] + e1[2][166] %3329;
                                                                                                                                                                                 u[2][167] = in_3[167] + e1[2][167] %3329;
                                                                                                                                                                                 u[2][168] = in_3[168] + e1[2][168] %3329;
                                                                                                                                                                                 u[2][169] = in_3[169] + e1[2][169] %3329;
                                                                                                                                                                                 u[2][170] = in_3[170] + e1[2][170] %3329;
                                                                                                                                                                                 u[2][171] = in_3[171] + e1[2][171] %3329;
                                                                                                                                                                                 u[2][172] = in_3[172] + e1[2][172] %3329;
                                                                                                                                                                                 u[2][173] = in_3[173] + e1[2][173] %3329;
                                                                                                                                                                                 u[2][174] = in_3[174] + e1[2][174] %3329;
                                                                                                                                                                                 u[2][175] = in_3[175] + e1[2][175] %3329;
                                                                                                                                                                                 u[2][176] = in_3[176] + e1[2][176] %3329;
                                                                                                                                                                                 u[2][177] = in_3[177] + e1[2][177] %3329;
                                                                                                                                                                                 u[2][178] = in_3[178] + e1[2][178] %3329;
                                                                                                                                                                                 u[2][179] = in_3[179] + e1[2][179] %3329;
                                                                                                                                                                                 u[2][180] = in_3[180] + e1[2][180] %3329;
                                                                                                                                                                                 u[2][181] = in_3[181] + e1[2][181] %3329;
                                                                                                                                                                                 u[2][182] = in_3[182] + e1[2][182] %3329;
                                                                                                                                                                                 u[2][183] = in_3[183] + e1[2][183] %3329;
                                                                                                                                                                                 u[2][184] = in_3[184] + e1[2][184] %3329;
                                                                                                                                                                                 u[2][185] = in_3[185] + e1[2][185] %3329;
                                                                                                                                                                                 u[2][186] = in_3[186] + e1[2][186] %3329;
                                                                                                                                                                                 u[2][187] = in_3[187] + e1[2][187] %3329;
                                                                                                                                                                                 u[2][188] = in_3[188] + e1[2][188] %3329;
                                                                                                                                                                                 u[2][189] = in_3[189] + e1[2][189] %3329;
                                                                                                                                                                                 u[2][190] = in_3[190] + e1[2][190] %3329;
                                                                                                                                                                                 u[2][191] = in_3[191] + e1[2][191] %3329;
                                                                                                                                                                                 u[2][192] = in_3[192] + e1[2][192] %3329;
                                                                                                                                                                                 u[2][193] = in_3[193] + e1[2][193] %3329;
                                                                                                                                                                                 u[2][194] = in_3[194] + e1[2][194] %3329;
                                                                                                                                                                                 u[2][195] = in_3[195] + e1[2][195] %3329;
                                                                                                                                                                                 u[2][196] = in_3[196] + e1[2][196] %3329;
                                                                                                                                                                                 u[2][197] = in_3[197] + e1[2][197] %3329;
                                                                                                                                                                                 u[2][198] = in_3[198] + e1[2][198] %3329;
                                                                                                                                                                                 u[2][199] = in_3[199] + e1[2][199] %3329;
                                                                                                                                                                                 u[2][200] = in_3[200] + e1[2][200] %3329;
                                                                                                                                                                                 u[2][201] = in_3[201] + e1[2][201] %3329;
                                                                                                                                                                                 u[2][202] = in_3[202] + e1[2][202] %3329;
                                                                                                                                                                                 u[2][203] = in_3[203] + e1[2][203] %3329;
                                                                                                                                                                                 u[2][204] = in_3[204] + e1[2][204] %3329;
                                                                                                                                                                                 u[2][205] = in_3[205] + e1[2][205] %3329;
                                                                                                                                                                                 u[2][206] = in_3[206] + e1[2][206] %3329;
                                                                                                                                                                                 u[2][207] = in_3[207] + e1[2][207] %3329;
                                                                                                                                                                                 u[2][208] = in_3[208] + e1[2][208] %3329;
                                                                                                                                                                                 u[2][209] = in_3[209] + e1[2][209] %3329;
                                                                                                                                                                                 u[2][210] = in_3[210] + e1[2][210] %3329;
                                                                                                                                                                                 u[2][211] = in_3[211] + e1[2][211] %3329;
                                                                                                                                                                                 u[2][212] = in_3[212] + e1[2][212] %3329;
                                                                                                                                                                                 u[2][213] = in_3[213] + e1[2][213] %3329;
                                                                                                                                                                                 u[2][214] = in_3[214] + e1[2][214] %3329;
                                                                                                                                                                                 u[2][215] = in_3[215] + e1[2][215] %3329;
                                                                                                                                                                                 u[2][216] = in_3[216] + e1[2][216] %3329;
                                                                                                                                                                                 u[2][217] = in_3[217] + e1[2][217] %3329;
                                                                                                                                                                                 u[2][218] = in_3[218] + e1[2][218] %3329;
                                                                                                                                                                                 u[2][219] = in_3[219] + e1[2][219] %3329;
                                                                                                                                                                                 u[2][220] = in_3[220] + e1[2][220] %3329;
                                                                                                                                                                                 u[2][221] = in_3[221] + e1[2][221] %3329;
                                                                                                                                                                                 u[2][222] = in_3[222] + e1[2][222] %3329;
                                                                                                                                                                                 u[2][223] = in_3[223] + e1[2][223] %3329;
                                                                                                                                                                                 u[2][224] = in_3[224] + e1[2][224] %3329;
                                                                                                                                                                                 u[2][225] = in_3[225] + e1[2][225] %3329;
                                                                                                                                                                                 u[2][226] = in_3[226] + e1[2][226] %3329;
                                                                                                                                                                                 u[2][227] = in_3[227] + e1[2][227] %3329;
                                                                                                                                                                                 u[2][228] = in_3[228] + e1[2][228] %3329;
                                                                                                                                                                                 u[2][229] = in_3[229] + e1[2][229] %3329;
                                                                                                                                                                                 u[2][230] = in_3[230] + e1[2][230] %3329;
                                                                                                                                                                                 u[2][231] = in_3[231] + e1[2][231] %3329;
                                                                                                                                                                                 u[2][232] = in_3[232] + e1[2][232] %3329;
                                                                                                                                                                                 u[2][233] = in_3[233] + e1[2][233] %3329;
                                                                                                                                                                                 u[2][234] = in_3[234] + e1[2][234] %3329;
                                                                                                                                                                                 u[2][235] = in_3[235] + e1[2][235] %3329;
                                                                                                                                                                                 u[2][236] = in_3[236] + e1[2][236] %3329;
                                                                                                                                                                                 u[2][237] = in_3[237] + e1[2][237] %3329;
                                                                                                                                                                                 u[2][238] = in_3[238] + e1[2][238] %3329;
                                                                                                                                                                                 u[2][239] = in_3[239] + e1[2][239] %3329;
                                                                                                                                                                                 u[2][240] = in_3[240] + e1[2][240] %3329;
                                                                                                                                                                                 u[2][241] = in_3[241] + e1[2][241] %3329;
                                                                                                                                                                                 u[2][242] = in_3[242] + e1[2][242] %3329;
                                                                                                                                                                                 u[2][243] = in_3[243] + e1[2][243] %3329;
                                                                                                                                                                                 u[2][244] = in_3[244] + e1[2][244] %3329;
                                                                                                                                                                                 u[2][245] = in_3[245] + e1[2][245] %3329;
                                                                                                                                                                                 u[2][246] = in_3[246] + e1[2][246] %3329;
                                                                                                                                                                                 u[2][247] = in_3[247] + e1[2][247] %3329;
                                                                                                                                                                                 u[2][248] = in_3[248] + e1[2][248] %3329;
                                                                                                                                                                                 u[2][249] = in_3[249] + e1[2][249] %3329;
                                                                                                                                                                                 u[2][250] = in_3[250] + e1[2][250] %3329;
                                                                                                                                                                                 u[2][251] = in_3[251] + e1[2][251] %3329;
                                                                                                                                                                                 u[2][252] = in_3[252] + e1[2][252] %3329;
                                                                                                                                                                                 u[2][253] = in_3[253] + e1[2][253] %3329;
                                                                                                                                                                                 u[2][254] = in_3[254] + e1[2][254] %3329;
                                                                                                                                                                                 u[2][255] = in_3[255] + e1[2][255] %3329;
                                                                                                                                                                                 result[0][0] = decom_out[0][0]+ mul_add_t[0][0] + {4'b0000, e2[0]}%3329;
                                                                                                                                                                                     result[0][1] = decom_out[0][1]+ mul_add_t[0][1] + {4'b0000, e2[1]}%3329;
                                                                                                                                                                                     result[0][2] = decom_out[0][2]+ mul_add_t[0][2] + {4'b0000, e2[2]}%3329;
                                                                                                                                                                                     result[0][3] = decom_out[0][3]+ mul_add_t[0][3] + {4'b0000, e2[3]}%3329;
                                                                                                                                                                                     result[0][4] = decom_out[0][4]+ mul_add_t[0][4] + {4'b0000, e2[4]}%3329;
                                                                                                                                                                                     result[0][5] = decom_out[0][5]+ mul_add_t[0][5] + {4'b0000, e2[5]}%3329;
                                                                                                                                                                                     result[0][6] = decom_out[0][6]+ mul_add_t[0][6] + {4'b0000, e2[6]}%3329;
                                                                                                                                                                                     result[0][7] = decom_out[0][7]+ mul_add_t[0][7] + {4'b0000, e2[7]}%3329;
                                                                                                                                                                                     result[0][8] = decom_out[0][8]+ mul_add_t[0][8] + {4'b0000, e2[8]}%3329;
                                                                                                                                                                                     result[0][9] = decom_out[0][9]+ mul_add_t[0][9] + {4'b0000, e2[9]}%3329;
                                                                                                                                                                                     result[0][10] = decom_out[0][10]+ mul_add_t[0][10] + {4'b0000, e2[10]}%3329;
                                                                                                                                                                                     result[0][11] = decom_out[0][11]+ mul_add_t[0][11] + {4'b0000, e2[11]}%3329;
                                                                                                                                                                                     result[0][12] = decom_out[0][12]+ mul_add_t[0][12] + {4'b0000, e2[12]}%3329;
                                                                                                                                                                                     result[0][13] = decom_out[0][13]+ mul_add_t[0][13] + {4'b0000, e2[13]}%3329;
                                                                                                                                                                                     result[0][14] = decom_out[0][14]+ mul_add_t[0][14] + {4'b0000, e2[14]}%3329;
                                                                                                                                                                                     result[0][15] = decom_out[0][15]+ mul_add_t[0][15] + {4'b0000, e2[15]}%3329;
                                                                                                                                                                                     result[0][16] = decom_out[0][16]+ mul_add_t[0][16] + {4'b0000, e2[16]}%3329;
                                                                                                                                                                                     result[0][17] = decom_out[0][17]+ mul_add_t[0][17] + {4'b0000, e2[17]}%3329;
                                                                                                                                                                                     result[0][18] = decom_out[0][18]+ mul_add_t[0][18] + {4'b0000, e2[18]}%3329;
                                                                                                                                                                                     result[0][19] = decom_out[0][19]+ mul_add_t[0][19] + {4'b0000, e2[19]}%3329;
                                                                                                                                                                                     result[0][20] = decom_out[0][20]+ mul_add_t[0][20] + {4'b0000, e2[20]}%3329;
                                                                                                                                                                                     result[0][21] = decom_out[0][21]+ mul_add_t[0][21] + {4'b0000, e2[21]}%3329;
                                                                                                                                                                                     result[0][22] = decom_out[0][22]+ mul_add_t[0][22] + {4'b0000, e2[22]}%3329;
                                                                                                                                                                                     result[0][23] = decom_out[0][23]+ mul_add_t[0][23] + {4'b0000, e2[23]}%3329;
                                                                                                                                                                                     result[0][24] = decom_out[0][24]+ mul_add_t[0][24] + {4'b0000, e2[24]}%3329;
                                                                                                                                                                                     result[0][25] = decom_out[0][25]+ mul_add_t[0][25] + {4'b0000, e2[25]}%3329;
                                                                                                                                                                                     result[0][26] = decom_out[0][26]+ mul_add_t[0][26] + {4'b0000, e2[26]}%3329;
                                                                                                                                                                                     result[0][27] = decom_out[0][27]+ mul_add_t[0][27] + {4'b0000, e2[27]}%3329;
                                                                                                                                                                                     result[0][28] = decom_out[0][28]+ mul_add_t[0][28] + {4'b0000, e2[28]}%3329;
                                                                                                                                                                                     result[0][29] = decom_out[0][29]+ mul_add_t[0][29] + {4'b0000, e2[29]}%3329;
                                                                                                                                                                                     result[0][30] = decom_out[0][30]+ mul_add_t[0][30] + {4'b0000, e2[30]}%3329;
                                                                                                                                                                                     result[0][31] = decom_out[0][31]+ mul_add_t[0][31] + {4'b0000, e2[31]}%3329;
                                                                                                                                                                                     result[0][32] = decom_out[0][32]+ mul_add_t[0][32] + {4'b0000, e2[32]}%3329;
                                                                                                                                                                                     result[0][33] = decom_out[0][33]+ mul_add_t[0][33] + {4'b0000, e2[33]}%3329;
                                                                                                                                                                                     result[0][34] = decom_out[0][34]+ mul_add_t[0][34] + {4'b0000, e2[34]}%3329;
                                                                                                                                                                                     result[0][35] = decom_out[0][35]+ mul_add_t[0][35] + {4'b0000, e2[35]}%3329;
                                                                                                                                                                                     result[0][36] = decom_out[0][36]+ mul_add_t[0][36] + {4'b0000, e2[36]}%3329;
                                                                                                                                                                                     result[0][37] = decom_out[0][37]+ mul_add_t[0][37] + {4'b0000, e2[37]}%3329;
                                                                                                                                                                                     result[0][38] = decom_out[0][38]+ mul_add_t[0][38] + {4'b0000, e2[38]}%3329;
                                                                                                                                                                                     result[0][39] = decom_out[0][39]+ mul_add_t[0][39] + {4'b0000, e2[39]}%3329;
                                                                                                                                                                                     result[0][40] = decom_out[0][40]+ mul_add_t[0][40] + {4'b0000, e2[40]}%3329;
                                                                                                                                                                                     result[0][41] = decom_out[0][41]+ mul_add_t[0][41] + {4'b0000, e2[41]}%3329;
                                                                                                                                                                                     result[0][42] = decom_out[0][42]+ mul_add_t[0][42] + {4'b0000, e2[42]}%3329;
                                                                                                                                                                                     result[0][43] = decom_out[0][43]+ mul_add_t[0][43] + {4'b0000, e2[43]}%3329;
                                                                                                                                                                                     result[0][44] = decom_out[0][44]+ mul_add_t[0][44] + {4'b0000, e2[44]}%3329;
                                                                                                                                                                                     result[0][45] = decom_out[0][45]+ mul_add_t[0][45] + {4'b0000, e2[45]}%3329;
                                                                                                                                                                                     result[0][46] = decom_out[0][46]+ mul_add_t[0][46] + {4'b0000, e2[46]}%3329;
                                                                                                                                                                                     result[0][47] = decom_out[0][47]+ mul_add_t[0][47] + {4'b0000, e2[47]}%3329;
                                                                                                                                                                                     result[0][48] = decom_out[0][48]+ mul_add_t[0][48] + {4'b0000, e2[48]}%3329;
                                                                                                                                                                                     result[0][49] = decom_out[0][49]+ mul_add_t[0][49] + {4'b0000, e2[49]}%3329;
                                                                                                                                                                                     result[0][50] = decom_out[0][50]+ mul_add_t[0][50] + {4'b0000, e2[50]}%3329;
                                                                                                                                                                                     result[0][51] = decom_out[0][51]+ mul_add_t[0][51] + {4'b0000, e2[51]}%3329;
                                                                                                                                                                                     result[0][52] = decom_out[0][52]+ mul_add_t[0][52] + {4'b0000, e2[52]}%3329;
                                                                                                                                                                                     result[0][53] = decom_out[0][53]+ mul_add_t[0][53] + {4'b0000, e2[53]}%3329;
                                                                                                                                                                                     result[0][54] = decom_out[0][54]+ mul_add_t[0][54] + {4'b0000, e2[54]}%3329;
                                                                                                                                                                                     result[0][55] = decom_out[0][55]+ mul_add_t[0][55] + {4'b0000, e2[55]}%3329;
                                                                                                                                                                                     result[0][56] = decom_out[0][56]+ mul_add_t[0][56] + {4'b0000, e2[56]}%3329;
                                                                                                                                                                                     result[0][57] = decom_out[0][57]+ mul_add_t[0][57] + {4'b0000, e2[57]}%3329;
                                                                                                                                                                                     result[0][58] = decom_out[0][58]+ mul_add_t[0][58] + {4'b0000, e2[58]}%3329;
                                                                                                                                                                                     result[0][59] = decom_out[0][59]+ mul_add_t[0][59] + {4'b0000, e2[59]}%3329;
                                                                                                                                                                                     result[0][60] = decom_out[0][60]+ mul_add_t[0][60] + {4'b0000, e2[60]}%3329;
                                                                                                                                                                                     result[0][61] = decom_out[0][61]+ mul_add_t[0][61] + {4'b0000, e2[61]}%3329;
                                                                                                                                                                                     result[0][62] = decom_out[0][62]+ mul_add_t[0][62] + {4'b0000, e2[62]}%3329;
                                                                                                                                                                                     result[0][63] = decom_out[0][63]+ mul_add_t[0][63] + {4'b0000, e2[63]}%3329;
                                                                                                                                                                                     result[0][64] = decom_out[0][64]+ mul_add_t[0][64] + {4'b0000, e2[64]}%3329;
                                                                                                                                                                                     result[0][65] = decom_out[0][65]+ mul_add_t[0][65] + {4'b0000, e2[65]}%3329;
                                                                                                                                                                                     result[0][66] = decom_out[0][66]+ mul_add_t[0][66] + {4'b0000, e2[66]}%3329;
                                                                                                                                                                                     result[0][67] = decom_out[0][67]+ mul_add_t[0][67] + {4'b0000, e2[67]}%3329;
                                                                                                                                                                                     result[0][68] = decom_out[0][68]+ mul_add_t[0][68] + {4'b0000, e2[68]}%3329;
                                                                                                                                                                                     result[0][69] = decom_out[0][69]+ mul_add_t[0][69] + {4'b0000, e2[69]}%3329;
                                                                                                                                                                                     result[0][70] = decom_out[0][70]+ mul_add_t[0][70] + {4'b0000, e2[70]}%3329;
                                                                                                                                                                                     result[0][71] = decom_out[0][71]+ mul_add_t[0][71] + {4'b0000, e2[71]}%3329;
                                                                                                                                                                                     result[0][72] = decom_out[0][72]+ mul_add_t[0][72] + {4'b0000, e2[72]}%3329;
                                                                                                                                                                                     result[0][73] = decom_out[0][73]+ mul_add_t[0][73] + {4'b0000, e2[73]}%3329;
                                                                                                                                                                                     result[0][74] = decom_out[0][74]+ mul_add_t[0][74] + {4'b0000, e2[74]}%3329;
                                                                                                                                                                                     result[0][75] = decom_out[0][75]+ mul_add_t[0][75] + {4'b0000, e2[75]}%3329;
                                                                                                                                                                                     result[0][76] = decom_out[0][76]+ mul_add_t[0][76] + {4'b0000, e2[76]}%3329;
                                                                                                                                                                                     result[0][77] = decom_out[0][77]+ mul_add_t[0][77] + {4'b0000, e2[77]}%3329;
                                                                                                                                                                                     result[0][78] = decom_out[0][78]+ mul_add_t[0][78] + {4'b0000, e2[78]}%3329;
                                                                                                                                                                                     result[0][79] = decom_out[0][79]+ mul_add_t[0][79] + {4'b0000, e2[79]}%3329;
                                                                                                                                                                                     result[0][80] = decom_out[0][80]+ mul_add_t[0][80] + {4'b0000, e2[80]}%3329;
                                                                                                                                                                                     result[0][81] = decom_out[0][81]+ mul_add_t[0][81] + {4'b0000, e2[81]}%3329;
                                                                                                                                                                                     result[0][82] = decom_out[0][82]+ mul_add_t[0][82] + {4'b0000, e2[82]}%3329;
                                                                                                                                                                                     result[0][83] = decom_out[0][83]+ mul_add_t[0][83] + {4'b0000, e2[83]}%3329;
                                                                                                                                                                                     result[0][84] = decom_out[0][84]+ mul_add_t[0][84] + {4'b0000, e2[84]}%3329;
                                                                                                                                                                                     result[0][85] = decom_out[0][85]+ mul_add_t[0][85] + {4'b0000, e2[85]}%3329;
                                                                                                                                                                                     result[0][86] = decom_out[0][86]+ mul_add_t[0][86] + {4'b0000, e2[86]}%3329;
                                                                                                                                                                                     result[0][87] = decom_out[0][87]+ mul_add_t[0][87] + {4'b0000, e2[87]}%3329;
                                                                                                                                                                                     result[0][88] = decom_out[0][88]+ mul_add_t[0][88] + {4'b0000, e2[88]}%3329;
                                                                                                                                                                                     result[0][89] = decom_out[0][89]+ mul_add_t[0][89] + {4'b0000, e2[89]}%3329;
                                                                                                                                                                                     result[0][90] = decom_out[0][90]+ mul_add_t[0][90] + {4'b0000, e2[90]}%3329;
                                                                                                                                                                                     result[0][91] = decom_out[0][91]+ mul_add_t[0][91] + {4'b0000, e2[91]}%3329;
                                                                                                                                                                                     result[0][92] = decom_out[0][92]+ mul_add_t[0][92] + {4'b0000, e2[92]}%3329;
                                                                                                                                                                                     result[0][93] = decom_out[0][93]+ mul_add_t[0][93] + {4'b0000, e2[93]}%3329;
                                                                                                                                                                                     result[0][94] = decom_out[0][94]+ mul_add_t[0][94] + {4'b0000, e2[94]}%3329;
                                                                                                                                                                                     result[0][95] = decom_out[0][95]+ mul_add_t[0][95] + {4'b0000, e2[95]}%3329;
                                                                                                                                                                                     result[0][96] = decom_out[0][96]+ mul_add_t[0][96] + {4'b0000, e2[96]}%3329;
                                                                                                                                                                                     result[0][97] = decom_out[0][97]+ mul_add_t[0][97] + {4'b0000, e2[97]}%3329;
                                                                                                                                                                                     result[0][98] = decom_out[0][98]+ mul_add_t[0][98] + {4'b0000, e2[98]}%3329;
                                                                                                                                                                                     result[0][99] = decom_out[0][99]+ mul_add_t[0][99] + {4'b0000, e2[99]}%3329;
                                                                                                                                                                                     result[0][100] = decom_out[0][100]+ mul_add_t[0][100] + {4'b0000, e2[100]}%3329;
                                                                                                                                                                                     result[0][101] = decom_out[0][101]+ mul_add_t[0][101] + {4'b0000, e2[101]}%3329;
                                                                                                                                                                                     result[0][102] = decom_out[0][102]+ mul_add_t[0][102] + {4'b0000, e2[102]}%3329;
                                                                                                                                                                                     result[0][103] = decom_out[0][103]+ mul_add_t[0][103] + {4'b0000, e2[103]}%3329;
                                                                                                                                                                                     result[0][104] = decom_out[0][104]+ mul_add_t[0][104] + {4'b0000, e2[104]}%3329;
                                                                                                                                                                                     result[0][105] = decom_out[0][105]+ mul_add_t[0][105] + {4'b0000, e2[105]}%3329;
                                                                                                                                                                                     result[0][106] = decom_out[0][106]+ mul_add_t[0][106] + {4'b0000, e2[106]}%3329;
                                                                                                                                                                                     result[0][107] = decom_out[0][107]+ mul_add_t[0][107] + {4'b0000, e2[107]}%3329;
                                                                                                                                                                                     result[0][108] = decom_out[0][108]+ mul_add_t[0][108] + {4'b0000, e2[108]}%3329;
                                                                                                                                                                                     result[0][109] = decom_out[0][109]+ mul_add_t[0][109] + {4'b0000, e2[109]}%3329;
                                                                                                                                                                                     result[0][110] = decom_out[0][110]+ mul_add_t[0][110] + {4'b0000, e2[110]}%3329;
                                                                                                                                                                                     result[0][111] = decom_out[0][111]+ mul_add_t[0][111] + {4'b0000, e2[111]}%3329;
                                                                                                                                                                                     result[0][112] = decom_out[0][112]+ mul_add_t[0][112] + {4'b0000, e2[112]}%3329;
                                                                                                                                                                                     result[0][113] = decom_out[0][113]+ mul_add_t[0][113] + {4'b0000, e2[113]}%3329;
                                                                                                                                                                                     result[0][114] = decom_out[0][114]+ mul_add_t[0][114] + {4'b0000, e2[114]}%3329;
                                                                                                                                                                                     result[0][115] = decom_out[0][115]+ mul_add_t[0][115] + {4'b0000, e2[115]}%3329;
                                                                                                                                                                                     result[0][116] = decom_out[0][116]+ mul_add_t[0][116] + {4'b0000, e2[116]}%3329;
                                                                                                                                                                                     result[0][117] = decom_out[0][117]+ mul_add_t[0][117] + {4'b0000, e2[117]}%3329;
                                                                                                                                                                                     result[0][118] = decom_out[0][118]+ mul_add_t[0][118] + {4'b0000, e2[118]}%3329;
                                                                                                                                                                                     result[0][119] = decom_out[0][119]+ mul_add_t[0][119] + {4'b0000, e2[119]}%3329;
                                                                                                                                                                                     result[0][120] = decom_out[0][120]+ mul_add_t[0][120] + {4'b0000, e2[120]}%3329;
                                                                                                                                                                                     result[0][121] = decom_out[0][121]+ mul_add_t[0][121] + {4'b0000, e2[121]}%3329;
                                                                                                                                                                                     result[0][122] = decom_out[0][122]+ mul_add_t[0][122] + {4'b0000, e2[122]}%3329;
                                                                                                                                                                                     result[0][123] = decom_out[0][123]+ mul_add_t[0][123] + {4'b0000, e2[123]}%3329;
                                                                                                                                                                                     result[0][124] = decom_out[0][124]+ mul_add_t[0][124] + {4'b0000, e2[124]}%3329;
                                                                                                                                                                                     result[0][125] = decom_out[0][125]+ mul_add_t[0][125] + {4'b0000, e2[125]}%3329;
                                                                                                                                                                                     result[0][126] = decom_out[0][126]+ mul_add_t[0][126] + {4'b0000, e2[126]}%3329;
                                                                                                                                                                                     result[0][127] = decom_out[0][127]+ mul_add_t[0][127] + {4'b0000, e2[127]}%3329;
                                                                                                                                                                                     result[0][128] = decom_out[0][128]+ mul_add_t[0][128] + {4'b0000, e2[128]}%3329;
                                                                                                                                                                                     result[0][129] = decom_out[0][129]+ mul_add_t[0][129] + {4'b0000, e2[129]}%3329;
                                                                                                                                                                                     result[0][130] = decom_out[0][130]+ mul_add_t[0][130] + {4'b0000, e2[130]}%3329;
                                                                                                                                                                                     result[0][131] = decom_out[0][131]+ mul_add_t[0][131] + {4'b0000, e2[131]}%3329;
                                                                                                                                                                                     result[0][132] = decom_out[0][132]+ mul_add_t[0][132] + {4'b0000, e2[132]}%3329;
                                                                                                                                                                                     result[0][133] = decom_out[0][133]+ mul_add_t[0][133] + {4'b0000, e2[133]}%3329;
                                                                                                                                                                                     result[0][134] = decom_out[0][134]+ mul_add_t[0][134] + {4'b0000, e2[134]}%3329;
                                                                                                                                                                                     result[0][135] = decom_out[0][135]+ mul_add_t[0][135] + {4'b0000, e2[135]}%3329;
                                                                                                                                                                                     result[0][136] = decom_out[0][136]+ mul_add_t[0][136] + {4'b0000, e2[136]}%3329;
                                                                                                                                                                                     result[0][137] = decom_out[0][137]+ mul_add_t[0][137] + {4'b0000, e2[137]}%3329;
                                                                                                                                                                                     result[0][138] = decom_out[0][138]+ mul_add_t[0][138] + {4'b0000, e2[138]}%3329;
                                                                                                                                                                                     result[0][139] = decom_out[0][139]+ mul_add_t[0][139] + {4'b0000, e2[139]}%3329;
                                                                                                                                                                                     result[0][140] = decom_out[0][140]+ mul_add_t[0][140] + {4'b0000, e2[140]}%3329;
                                                                                                                                                                                     result[0][141] = decom_out[0][141]+ mul_add_t[0][141] + {4'b0000, e2[141]}%3329;
                                                                                                                                                                                     result[0][142] = decom_out[0][142]+ mul_add_t[0][142] + {4'b0000, e2[142]}%3329;
                                                                                                                                                                                     result[0][143] = decom_out[0][143]+ mul_add_t[0][143] + {4'b0000, e2[143]}%3329;
                                                                                                                                                                                     result[0][144] = decom_out[0][144]+ mul_add_t[0][144] + {4'b0000, e2[144]}%3329;
                                                                                                                                                                                     result[0][145] = decom_out[0][145]+ mul_add_t[0][145] + {4'b0000, e2[145]}%3329;
                                                                                                                                                                                     result[0][146] = decom_out[0][146]+ mul_add_t[0][146] + {4'b0000, e2[146]}%3329;
                                                                                                                                                                                     result[0][147] = decom_out[0][147]+ mul_add_t[0][147] + {4'b0000, e2[147]}%3329;
                                                                                                                                                                                     result[0][148] = decom_out[0][148]+ mul_add_t[0][148] + {4'b0000, e2[148]}%3329;
                                                                                                                                                                                     result[0][149] = decom_out[0][149]+ mul_add_t[0][149] + {4'b0000, e2[149]}%3329;
                                                                                                                                                                                     result[0][150] = decom_out[0][150]+ mul_add_t[0][150] + {4'b0000, e2[150]}%3329;
                                                                                                                                                                                     result[0][151] = decom_out[0][151]+ mul_add_t[0][151] + {4'b0000, e2[151]}%3329;
                                                                                                                                                                                     result[0][152] = decom_out[0][152]+ mul_add_t[0][152] + {4'b0000, e2[152]}%3329;
                                                                                                                                                                                     result[0][153] = decom_out[0][153]+ mul_add_t[0][153] + {4'b0000, e2[153]}%3329;
                                                                                                                                                                                     result[0][154] = decom_out[0][154]+ mul_add_t[0][154] + {4'b0000, e2[154]}%3329;
                                                                                                                                                                                     result[0][155] = decom_out[0][155]+ mul_add_t[0][155] + {4'b0000, e2[155]}%3329;
                                                                                                                                                                                     result[0][156] = decom_out[0][156]+ mul_add_t[0][156] + {4'b0000, e2[156]}%3329;
                                                                                                                                                                                     result[0][157] = decom_out[0][157]+ mul_add_t[0][157] + {4'b0000, e2[157]}%3329;
                                                                                                                                                                                     result[0][158] = decom_out[0][158]+ mul_add_t[0][158] + {4'b0000, e2[158]}%3329;
                                                                                                                                                                                     result[0][159] = decom_out[0][159]+ mul_add_t[0][159] + {4'b0000, e2[159]}%3329;
                                                                                                                                                                                     result[0][160] = decom_out[0][160]+ mul_add_t[0][160] + {4'b0000, e2[160]}%3329;
                                                                                                                                                                                     result[0][161] = decom_out[0][161]+ mul_add_t[0][161] + {4'b0000, e2[161]}%3329;
                                                                                                                                                                                     result[0][162] = decom_out[0][162]+ mul_add_t[0][162] + {4'b0000, e2[162]}%3329;
                                                                                                                                                                                     result[0][163] = decom_out[0][163]+ mul_add_t[0][163] + {4'b0000, e2[163]}%3329;
                                                                                                                                                                                     result[0][164] = decom_out[0][164]+ mul_add_t[0][164] + {4'b0000, e2[164]}%3329;
                                                                                                                                                                                     result[0][165] = decom_out[0][165]+ mul_add_t[0][165] + {4'b0000, e2[165]}%3329;
                                                                                                                                                                                     result[0][166] = decom_out[0][166]+ mul_add_t[0][166] + {4'b0000, e2[166]}%3329;
                                                                                                                                                                                     result[0][167] = decom_out[0][167]+ mul_add_t[0][167] + {4'b0000, e2[167]}%3329;
                                                                                                                                                                                     result[0][168] = decom_out[0][168]+ mul_add_t[0][168] + {4'b0000, e2[168]}%3329;
                                                                                                                                                                                     result[0][169] = decom_out[0][169]+ mul_add_t[0][169] + {4'b0000, e2[169]}%3329;
                                                                                                                                                                                     result[0][170] = decom_out[0][170]+ mul_add_t[0][170] + {4'b0000, e2[170]}%3329;
                                                                                                                                                                                     result[0][171] = decom_out[0][171]+ mul_add_t[0][171] + {4'b0000, e2[171]}%3329;
                                                                                                                                                                                     result[0][172] = decom_out[0][172]+ mul_add_t[0][172] + {4'b0000, e2[172]}%3329;
                                                                                                                                                                                     result[0][173] = decom_out[0][173]+ mul_add_t[0][173] + {4'b0000, e2[173]}%3329;
                                                                                                                                                                                     result[0][174] = decom_out[0][174]+ mul_add_t[0][174] + {4'b0000, e2[174]}%3329;
                                                                                                                                                                                     result[0][175] = decom_out[0][175]+ mul_add_t[0][175] + {4'b0000, e2[175]}%3329;
                                                                                                                                                                                     result[0][176] = decom_out[0][176]+ mul_add_t[0][176] + {4'b0000, e2[176]}%3329;
                                                                                                                                                                                     result[0][177] = decom_out[0][177]+ mul_add_t[0][177] + {4'b0000, e2[177]}%3329;
                                                                                                                                                                                     result[0][178] = decom_out[0][178]+ mul_add_t[0][178] + {4'b0000, e2[178]}%3329;
                                                                                                                                                                                     result[0][179] = decom_out[0][179]+ mul_add_t[0][179] + {4'b0000, e2[179]}%3329;
                                                                                                                                                                                     result[0][180] = decom_out[0][180]+ mul_add_t[0][180] + {4'b0000, e2[180]}%3329;
                                                                                                                                                                                     result[0][181] = decom_out[0][181]+ mul_add_t[0][181] + {4'b0000, e2[181]}%3329;
                                                                                                                                                                                     result[0][182] = decom_out[0][182]+ mul_add_t[0][182] + {4'b0000, e2[182]}%3329;
                                                                                                                                                                                     result[0][183] = decom_out[0][183]+ mul_add_t[0][183] + {4'b0000, e2[183]}%3329;
                                                                                                                                                                                     result[0][184] = decom_out[0][184]+ mul_add_t[0][184] + {4'b0000, e2[184]}%3329;
                                                                                                                                                                                     result[0][185] = decom_out[0][185]+ mul_add_t[0][185] + {4'b0000, e2[185]}%3329;
                                                                                                                                                                                     result[0][186] = decom_out[0][186]+ mul_add_t[0][186] + {4'b0000, e2[186]}%3329;
                                                                                                                                                                                     result[0][187] = decom_out[0][187]+ mul_add_t[0][187] + {4'b0000, e2[187]}%3329;
                                                                                                                                                                                     result[0][188] = decom_out[0][188]+ mul_add_t[0][188] + {4'b0000, e2[188]}%3329;
                                                                                                                                                                                     result[0][189] = decom_out[0][189]+ mul_add_t[0][189] + {4'b0000, e2[189]}%3329;
                                                                                                                                                                                     result[0][190] = decom_out[0][190]+ mul_add_t[0][190] + {4'b0000, e2[190]}%3329;
                                                                                                                                                                                     result[0][191] = decom_out[0][191]+ mul_add_t[0][191] + {4'b0000, e2[191]}%3329;
                                                                                                                                                                                     result[0][192] = decom_out[0][192]+ mul_add_t[0][192] + {4'b0000, e2[192]}%3329;
                                                                                                                                                                                     result[0][193] = decom_out[0][193]+ mul_add_t[0][193] + {4'b0000, e2[193]}%3329;
                                                                                                                                                                                     result[0][194] = decom_out[0][194]+ mul_add_t[0][194] + {4'b0000, e2[194]}%3329;
                                                                                                                                                                                     result[0][195] = decom_out[0][195]+ mul_add_t[0][195] + {4'b0000, e2[195]}%3329;
                                                                                                                                                                                     result[0][196] = decom_out[0][196]+ mul_add_t[0][196] + {4'b0000, e2[196]}%3329;
                                                                                                                                                                                     result[0][197] = decom_out[0][197]+ mul_add_t[0][197] + {4'b0000, e2[197]}%3329;
                                                                                                                                                                                     result[0][198] = decom_out[0][198]+ mul_add_t[0][198] + {4'b0000, e2[198]}%3329;
                                                                                                                                                                                     result[0][199] = decom_out[0][199]+ mul_add_t[0][199] + {4'b0000, e2[199]}%3329;
                                                                                                                                                                                     result[0][200] = decom_out[0][200]+ mul_add_t[0][200] + {4'b0000, e2[200]}%3329;
                                                                                                                                                                                     result[0][201] = decom_out[0][201]+ mul_add_t[0][201] + {4'b0000, e2[201]}%3329;
                                                                                                                                                                                     result[0][202] = decom_out[0][202]+ mul_add_t[0][202] + {4'b0000, e2[202]}%3329;
                                                                                                                                                                                     result[0][203] = decom_out[0][203]+ mul_add_t[0][203] + {4'b0000, e2[203]}%3329;
                                                                                                                                                                                     result[0][204] = decom_out[0][204]+ mul_add_t[0][204] + {4'b0000, e2[204]}%3329;
                                                                                                                                                                                     result[0][205] = decom_out[0][205]+ mul_add_t[0][205] + {4'b0000, e2[205]}%3329;
                                                                                                                                                                                     result[0][206] = decom_out[0][206]+ mul_add_t[0][206] + {4'b0000, e2[206]}%3329;
                                                                                                                                                                                     result[0][207] = decom_out[0][207]+ mul_add_t[0][207] + {4'b0000, e2[207]}%3329;
                                                                                                                                                                                     result[0][208] = decom_out[0][208]+ mul_add_t[0][208] + {4'b0000, e2[208]}%3329;
                                                                                                                                                                                     result[0][209] = decom_out[0][209]+ mul_add_t[0][209] + {4'b0000, e2[209]}%3329;
                                                                                                                                                                                     result[0][210] = decom_out[0][210]+ mul_add_t[0][210] + {4'b0000, e2[210]}%3329;
                                                                                                                                                                                     result[0][211] = decom_out[0][211]+ mul_add_t[0][211] + {4'b0000, e2[211]}%3329;
                                                                                                                                                                                     result[0][212] = decom_out[0][212]+ mul_add_t[0][212] + {4'b0000, e2[212]}%3329;
                                                                                                                                                                                     result[0][213] = decom_out[0][213]+ mul_add_t[0][213] + {4'b0000, e2[213]}%3329;
                                                                                                                                                                                     result[0][214] = decom_out[0][214]+ mul_add_t[0][214] + {4'b0000, e2[214]}%3329;
                                                                                                                                                                                     result[0][215] = decom_out[0][215]+ mul_add_t[0][215] + {4'b0000, e2[215]}%3329;
                                                                                                                                                                                     result[0][216] = decom_out[0][216]+ mul_add_t[0][216] + {4'b0000, e2[216]}%3329;
                                                                                                                                                                                     result[0][217] = decom_out[0][217]+ mul_add_t[0][217] + {4'b0000, e2[217]}%3329;
                                                                                                                                                                                     result[0][218] = decom_out[0][218]+ mul_add_t[0][218] + {4'b0000, e2[218]}%3329;
                                                                                                                                                                                     result[0][219] = decom_out[0][219]+ mul_add_t[0][219] + {4'b0000, e2[219]}%3329;
                                                                                                                                                                                     result[0][220] = decom_out[0][220]+ mul_add_t[0][220] + {4'b0000, e2[220]}%3329;
                                                                                                                                                                                     result[0][221] = decom_out[0][221]+ mul_add_t[0][221] + {4'b0000, e2[221]}%3329;
                                                                                                                                                                                     result[0][222] = decom_out[0][222]+ mul_add_t[0][222] + {4'b0000, e2[222]}%3329;
                                                                                                                                                                                     result[0][223] = decom_out[0][223]+ mul_add_t[0][223] + {4'b0000, e2[223]}%3329;
                                                                                                                                                                                     result[0][224] = decom_out[0][224]+ mul_add_t[0][224] + {4'b0000, e2[224]}%3329;
                                                                                                                                                                                     result[0][225] = decom_out[0][225]+ mul_add_t[0][225] + {4'b0000, e2[225]}%3329;
                                                                                                                                                                                     result[0][226] = decom_out[0][226]+ mul_add_t[0][226] + {4'b0000, e2[226]}%3329;
                                                                                                                                                                                     result[0][227] = decom_out[0][227]+ mul_add_t[0][227] + {4'b0000, e2[227]}%3329;
                                                                                                                                                                                     result[0][228] = decom_out[0][228]+ mul_add_t[0][228] + {4'b0000, e2[228]}%3329;
                                                                                                                                                                                     result[0][229] = decom_out[0][229]+ mul_add_t[0][229] + {4'b0000, e2[229]}%3329;
                                                                                                                                                                                     result[0][230] = decom_out[0][230]+ mul_add_t[0][230] + {4'b0000, e2[230]}%3329;
                                                                                                                                                                                     result[0][231] = decom_out[0][231]+ mul_add_t[0][231] + {4'b0000, e2[231]}%3329;
                                                                                                                                                                                     result[0][232] = decom_out[0][232]+ mul_add_t[0][232] + {4'b0000, e2[232]}%3329;
                                                                                                                                                                                     result[0][233] = decom_out[0][233]+ mul_add_t[0][233] + {4'b0000, e2[233]}%3329;
                                                                                                                                                                                     result[0][234] = decom_out[0][234]+ mul_add_t[0][234] + {4'b0000, e2[234]}%3329;
                                                                                                                                                                                     result[0][235] = decom_out[0][235]+ mul_add_t[0][235] + {4'b0000, e2[235]}%3329;
                                                                                                                                                                                     result[0][236] = decom_out[0][236]+ mul_add_t[0][236] + {4'b0000, e2[236]}%3329;
                                                                                                                                                                                     result[0][237] = decom_out[0][237]+ mul_add_t[0][237] + {4'b0000, e2[237]}%3329;
                                                                                                                                                                                     result[0][238] = decom_out[0][238]+ mul_add_t[0][238] + {4'b0000, e2[238]}%3329;
                                                                                                                                                                                     result[0][239] = decom_out[0][239]+ mul_add_t[0][239] + {4'b0000, e2[239]}%3329;
                                                                                                                                                                                     result[0][240] = decom_out[0][240]+ mul_add_t[0][240] + {4'b0000, e2[240]}%3329;
                                                                                                                                                                                     result[0][241] = decom_out[0][241]+ mul_add_t[0][241] + {4'b0000, e2[241]}%3329;
                                                                                                                                                                                     result[0][242] = decom_out[0][242]+ mul_add_t[0][242] + {4'b0000, e2[242]}%3329;
                                                                                                                                                                                     result[0][243] = decom_out[0][243]+ mul_add_t[0][243] + {4'b0000, e2[243]}%3329;
                                                                                                                                                                                     result[0][244] = decom_out[0][244]+ mul_add_t[0][244] + {4'b0000, e2[244]}%3329;
                                                                                                                                                                                     result[0][245] = decom_out[0][245]+ mul_add_t[0][245] + {4'b0000, e2[245]}%3329;
                                                                                                                                                                                     result[0][246] = decom_out[0][246]+ mul_add_t[0][246] + {4'b0000, e2[246]}%3329;
                                                                                                                                                                                     result[0][247] = decom_out[0][247]+ mul_add_t[0][247] + {4'b0000, e2[247]}%3329;
                                                                                                                                                                                     result[0][248] = decom_out[0][248]+ mul_add_t[0][248] + {4'b0000, e2[248]}%3329;
                                                                                                                                                                                     result[0][249] = decom_out[0][249]+ mul_add_t[0][249] + {4'b0000, e2[249]}%3329;
                                                                                                                                                                                     result[0][250] = decom_out[0][250]+ mul_add_t[0][250] + {4'b0000, e2[250]}%3329;
                                                                                                                                                                                     result[0][251] = decom_out[0][251]+ mul_add_t[0][251] + {4'b0000, e2[251]}%3329;
                                                                                                                                                                                     result[0][252] = decom_out[0][252]+ mul_add_t[0][252] + {4'b0000, e2[252]}%3329;
                                                                                                                                                                                     result[0][253] = decom_out[0][253]+ mul_add_t[0][253] + {4'b0000, e2[253]}%3329;
                                                                                                                                                                                     result[0][254] = decom_out[0][254]+ mul_add_t[0][254] + {4'b0000, e2[254]}%3329;
                                                                                                                                                                                     result[0][255] = decom_out[0][255]+ mul_add_t[0][255] + {4'b0000, e2[255]}%3329;
                                                                                                                                                                                     result[1][0] = decom_out[1][0]+ mul_add_t[1][0] + {4'b0000, e2[0]}%3329;
                                                                                                                                                                                     result[1][1] = decom_out[1][1]+ mul_add_t[1][1] + {4'b0000, e2[1]}%3329;
                                                                                                                                                                                     result[1][2] = decom_out[1][2]+ mul_add_t[1][2] + {4'b0000, e2[2]}%3329;
                                                                                                                                                                                     result[1][3] = decom_out[1][3]+ mul_add_t[1][3] + {4'b0000, e2[3]}%3329;
                                                                                                                                                                                     result[1][4] = decom_out[1][4]+ mul_add_t[1][4] + {4'b0000, e2[4]}%3329;
                                                                                                                                                                                     result[1][5] = decom_out[1][5]+ mul_add_t[1][5] + {4'b0000, e2[5]}%3329;
                                                                                                                                                                                     result[1][6] = decom_out[1][6]+ mul_add_t[1][6] + {4'b0000, e2[6]}%3329;
                                                                                                                                                                                     result[1][7] = decom_out[1][7]+ mul_add_t[1][7] + {4'b0000, e2[7]}%3329;
                                                                                                                                                                                     result[1][8] = decom_out[1][8]+ mul_add_t[1][8] + {4'b0000, e2[8]}%3329;
                                                                                                                                                                                     result[1][9] = decom_out[1][9]+ mul_add_t[1][9] + {4'b0000, e2[9]}%3329;
                                                                                                                                                                                     result[1][10] = decom_out[1][10]+ mul_add_t[1][10] + {4'b0000, e2[10]}%3329;
                                                                                                                                                                                     result[1][11] = decom_out[1][11]+ mul_add_t[1][11] + {4'b0000, e2[11]}%3329;
                                                                                                                                                                                     result[1][12] = decom_out[1][12]+ mul_add_t[1][12] + {4'b0000, e2[12]}%3329;
                                                                                                                                                                                     result[1][13] = decom_out[1][13]+ mul_add_t[1][13] + {4'b0000, e2[13]}%3329;
                                                                                                                                                                                     result[1][14] = decom_out[1][14]+ mul_add_t[1][14] + {4'b0000, e2[14]}%3329;
                                                                                                                                                                                     result[1][15] = decom_out[1][15]+ mul_add_t[1][15] + {4'b0000, e2[15]}%3329;
                                                                                                                                                                                     result[1][16] = decom_out[1][16]+ mul_add_t[1][16] + {4'b0000, e2[16]}%3329;
                                                                                                                                                                                     result[1][17] = decom_out[1][17]+ mul_add_t[1][17] + {4'b0000, e2[17]}%3329;
                                                                                                                                                                                     result[1][18] = decom_out[1][18]+ mul_add_t[1][18] + {4'b0000, e2[18]}%3329;
                                                                                                                                                                                     result[1][19] = decom_out[1][19]+ mul_add_t[1][19] + {4'b0000, e2[19]}%3329;
                                                                                                                                                                                     result[1][20] = decom_out[1][20]+ mul_add_t[1][20] + {4'b0000, e2[20]}%3329;
                                                                                                                                                                                     result[1][21] = decom_out[1][21]+ mul_add_t[1][21] + {4'b0000, e2[21]}%3329;
                                                                                                                                                                                     result[1][22] = decom_out[1][22]+ mul_add_t[1][22] + {4'b0000, e2[22]}%3329;
                                                                                                                                                                                     result[1][23] = decom_out[1][23]+ mul_add_t[1][23] + {4'b0000, e2[23]}%3329;
                                                                                                                                                                                     result[1][24] = decom_out[1][24]+ mul_add_t[1][24] + {4'b0000, e2[24]}%3329;
                                                                                                                                                                                     result[1][25] = decom_out[1][25]+ mul_add_t[1][25] + {4'b0000, e2[25]}%3329;
                                                                                                                                                                                     result[1][26] = decom_out[1][26]+ mul_add_t[1][26] + {4'b0000, e2[26]}%3329;
                                                                                                                                                                                     result[1][27] = decom_out[1][27]+ mul_add_t[1][27] + {4'b0000, e2[27]}%3329;
                                                                                                                                                                                     result[1][28] = decom_out[1][28]+ mul_add_t[1][28] + {4'b0000, e2[28]}%3329;
                                                                                                                                                                                     result[1][29] = decom_out[1][29]+ mul_add_t[1][29] + {4'b0000, e2[29]}%3329;
                                                                                                                                                                                     result[1][30] = decom_out[1][30]+ mul_add_t[1][30] + {4'b0000, e2[30]}%3329;
                                                                                                                                                                                     result[1][31] = decom_out[1][31]+ mul_add_t[1][31] + {4'b0000, e2[31]}%3329;
                                                                                                                                                                                     result[1][32] = decom_out[1][32]+ mul_add_t[1][32] + {4'b0000, e2[32]}%3329;
                                                                                                                                                                                     result[1][33] = decom_out[1][33]+ mul_add_t[1][33] + {4'b0000, e2[33]}%3329;
                                                                                                                                                                                     result[1][34] = decom_out[1][34]+ mul_add_t[1][34] + {4'b0000, e2[34]}%3329;
                                                                                                                                                                                     result[1][35] = decom_out[1][35]+ mul_add_t[1][35] + {4'b0000, e2[35]}%3329;
                                                                                                                                                                                     result[1][36] = decom_out[1][36]+ mul_add_t[1][36] + {4'b0000, e2[36]}%3329;
                                                                                                                                                                                     result[1][37] = decom_out[1][37]+ mul_add_t[1][37] + {4'b0000, e2[37]}%3329;
                                                                                                                                                                                     result[1][38] = decom_out[1][38]+ mul_add_t[1][38] + {4'b0000, e2[38]}%3329;
                                                                                                                                                                                     result[1][39] = decom_out[1][39]+ mul_add_t[1][39] + {4'b0000, e2[39]}%3329;
                                                                                                                                                                                     result[1][40] = decom_out[1][40]+ mul_add_t[1][40] + {4'b0000, e2[40]}%3329;
                                                                                                                                                                                     result[1][41] = decom_out[1][41]+ mul_add_t[1][41] + {4'b0000, e2[41]}%3329;
                                                                                                                                                                                     result[1][42] = decom_out[1][42]+ mul_add_t[1][42] + {4'b0000, e2[42]}%3329;
                                                                                                                                                                                     result[1][43] = decom_out[1][43]+ mul_add_t[1][43] + {4'b0000, e2[43]}%3329;
                                                                                                                                                                                     result[1][44] = decom_out[1][44]+ mul_add_t[1][44] + {4'b0000, e2[44]}%3329;
                                                                                                                                                                                     result[1][45] = decom_out[1][45]+ mul_add_t[1][45] + {4'b0000, e2[45]}%3329;
                                                                                                                                                                                     result[1][46] = decom_out[1][46]+ mul_add_t[1][46] + {4'b0000, e2[46]}%3329;
                                                                                                                                                                                     result[1][47] = decom_out[1][47]+ mul_add_t[1][47] + {4'b0000, e2[47]}%3329;
                                                                                                                                                                                     result[1][48] = decom_out[1][48]+ mul_add_t[1][48] + {4'b0000, e2[48]}%3329;
                                                                                                                                                                                     result[1][49] = decom_out[1][49]+ mul_add_t[1][49] + {4'b0000, e2[49]}%3329;
                                                                                                                                                                                     result[1][50] = decom_out[1][50]+ mul_add_t[1][50] + {4'b0000, e2[50]}%3329;
                                                                                                                                                                                     result[1][51] = decom_out[1][51]+ mul_add_t[1][51] + {4'b0000, e2[51]}%3329;
                                                                                                                                                                                     result[1][52] = decom_out[1][52]+ mul_add_t[1][52] + {4'b0000, e2[52]}%3329;
                                                                                                                                                                                     result[1][53] = decom_out[1][53]+ mul_add_t[1][53] + {4'b0000, e2[53]}%3329;
                                                                                                                                                                                     result[1][54] = decom_out[1][54]+ mul_add_t[1][54] + {4'b0000, e2[54]}%3329;
                                                                                                                                                                                     result[1][55] = decom_out[1][55]+ mul_add_t[1][55] + {4'b0000, e2[55]}%3329;
                                                                                                                                                                                     result[1][56] = decom_out[1][56]+ mul_add_t[1][56] + {4'b0000, e2[56]}%3329;
                                                                                                                                                                                     result[1][57] = decom_out[1][57]+ mul_add_t[1][57] + {4'b0000, e2[57]}%3329;
                                                                                                                                                                                     result[1][58] = decom_out[1][58]+ mul_add_t[1][58] + {4'b0000, e2[58]}%3329;
                                                                                                                                                                                     result[1][59] = decom_out[1][59]+ mul_add_t[1][59] + {4'b0000, e2[59]}%3329;
                                                                                                                                                                                     result[1][60] = decom_out[1][60]+ mul_add_t[1][60] + {4'b0000, e2[60]}%3329;
                                                                                                                                                                                     result[1][61] = decom_out[1][61]+ mul_add_t[1][61] + {4'b0000, e2[61]}%3329;
                                                                                                                                                                                     result[1][62] = decom_out[1][62]+ mul_add_t[1][62] + {4'b0000, e2[62]}%3329;
                                                                                                                                                                                     result[1][63] = decom_out[1][63]+ mul_add_t[1][63] + {4'b0000, e2[63]}%3329;
                                                                                                                                                                                     result[1][64] = decom_out[1][64]+ mul_add_t[1][64] + {4'b0000, e2[64]}%3329;
                                                                                                                                                                                     result[1][65] = decom_out[1][65]+ mul_add_t[1][65] + {4'b0000, e2[65]}%3329;
                                                                                                                                                                                     result[1][66] = decom_out[1][66]+ mul_add_t[1][66] + {4'b0000, e2[66]}%3329;
                                                                                                                                                                                     result[1][67] = decom_out[1][67]+ mul_add_t[1][67] + {4'b0000, e2[67]}%3329;
                                                                                                                                                                                     result[1][68] = decom_out[1][68]+ mul_add_t[1][68] + {4'b0000, e2[68]}%3329;
                                                                                                                                                                                     result[1][69] = decom_out[1][69]+ mul_add_t[1][69] + {4'b0000, e2[69]}%3329;
                                                                                                                                                                                     result[1][70] = decom_out[1][70]+ mul_add_t[1][70] + {4'b0000, e2[70]}%3329;
                                                                                                                                                                                     result[1][71] = decom_out[1][71]+ mul_add_t[1][71] + {4'b0000, e2[71]}%3329;
                                                                                                                                                                                     result[1][72] = decom_out[1][72]+ mul_add_t[1][72] + {4'b0000, e2[72]}%3329;
                                                                                                                                                                                     result[1][73] = decom_out[1][73]+ mul_add_t[1][73] + {4'b0000, e2[73]}%3329;
                                                                                                                                                                                     result[1][74] = decom_out[1][74]+ mul_add_t[1][74] + {4'b0000, e2[74]}%3329;
                                                                                                                                                                                     result[1][75] = decom_out[1][75]+ mul_add_t[1][75] + {4'b0000, e2[75]}%3329;
                                                                                                                                                                                     result[1][76] = decom_out[1][76]+ mul_add_t[1][76] + {4'b0000, e2[76]}%3329;
                                                                                                                                                                                     result[1][77] = decom_out[1][77]+ mul_add_t[1][77] + {4'b0000, e2[77]}%3329;
                                                                                                                                                                                     result[1][78] = decom_out[1][78]+ mul_add_t[1][78] + {4'b0000, e2[78]}%3329;
                                                                                                                                                                                     result[1][79] = decom_out[1][79]+ mul_add_t[1][79] + {4'b0000, e2[79]}%3329;
                                                                                                                                                                                     result[1][80] = decom_out[1][80]+ mul_add_t[1][80] + {4'b0000, e2[80]}%3329;
                                                                                                                                                                                     result[1][81] = decom_out[1][81]+ mul_add_t[1][81] + {4'b0000, e2[81]}%3329;
                                                                                                                                                                                     result[1][82] = decom_out[1][82]+ mul_add_t[1][82] + {4'b0000, e2[82]}%3329;
                                                                                                                                                                                     result[1][83] = decom_out[1][83]+ mul_add_t[1][83] + {4'b0000, e2[83]}%3329;
                                                                                                                                                                                     result[1][84] = decom_out[1][84]+ mul_add_t[1][84] + {4'b0000, e2[84]}%3329;
                                                                                                                                                                                     result[1][85] = decom_out[1][85]+ mul_add_t[1][85] + {4'b0000, e2[85]}%3329;
                                                                                                                                                                                     result[1][86] = decom_out[1][86]+ mul_add_t[1][86] + {4'b0000, e2[86]}%3329;
                                                                                                                                                                                     result[1][87] = decom_out[1][87]+ mul_add_t[1][87] + {4'b0000, e2[87]}%3329;
                                                                                                                                                                                     result[1][88] = decom_out[1][88]+ mul_add_t[1][88] + {4'b0000, e2[88]}%3329;
                                                                                                                                                                                     result[1][89] = decom_out[1][89]+ mul_add_t[1][89] + {4'b0000, e2[89]}%3329;
                                                                                                                                                                                     result[1][90] = decom_out[1][90]+ mul_add_t[1][90] + {4'b0000, e2[90]}%3329;
                                                                                                                                                                                     result[1][91] = decom_out[1][91]+ mul_add_t[1][91] + {4'b0000, e2[91]}%3329;
                                                                                                                                                                                     result[1][92] = decom_out[1][92]+ mul_add_t[1][92] + {4'b0000, e2[92]}%3329;
                                                                                                                                                                                     result[1][93] = decom_out[1][93]+ mul_add_t[1][93] + {4'b0000, e2[93]}%3329;
                                                                                                                                                                                     result[1][94] = decom_out[1][94]+ mul_add_t[1][94] + {4'b0000, e2[94]}%3329;
                                                                                                                                                                                     result[1][95] = decom_out[1][95]+ mul_add_t[1][95] + {4'b0000, e2[95]}%3329;
                                                                                                                                                                                     result[1][96] = decom_out[1][96]+ mul_add_t[1][96] + {4'b0000, e2[96]}%3329;
                                                                                                                                                                                     result[1][97] = decom_out[1][97]+ mul_add_t[1][97] + {4'b0000, e2[97]}%3329;
                                                                                                                                                                                     result[1][98] = decom_out[1][98]+ mul_add_t[1][98] + {4'b0000, e2[98]}%3329;
                                                                                                                                                                                     result[1][99] = decom_out[1][99]+ mul_add_t[1][99] + {4'b0000, e2[99]}%3329;
                                                                                                                                                                                     result[1][100] = decom_out[1][100]+ mul_add_t[1][100] + {4'b0000, e2[100]}%3329;
                                                                                                                                                                                     result[1][101] = decom_out[1][101]+ mul_add_t[1][101] + {4'b0000, e2[101]}%3329;
                                                                                                                                                                                     result[1][102] = decom_out[1][102]+ mul_add_t[1][102] + {4'b0000, e2[102]}%3329;
                                                                                                                                                                                     result[1][103] = decom_out[1][103]+ mul_add_t[1][103] + {4'b0000, e2[103]}%3329;
                                                                                                                                                                                     result[1][104] = decom_out[1][104]+ mul_add_t[1][104] + {4'b0000, e2[104]}%3329;
                                                                                                                                                                                     result[1][105] = decom_out[1][105]+ mul_add_t[1][105] + {4'b0000, e2[105]}%3329;
                                                                                                                                                                                     result[1][106] = decom_out[1][106]+ mul_add_t[1][106] + {4'b0000, e2[106]}%3329;
                                                                                                                                                                                     result[1][107] = decom_out[1][107]+ mul_add_t[1][107] + {4'b0000, e2[107]}%3329;
                                                                                                                                                                                     result[1][108] = decom_out[1][108]+ mul_add_t[1][108] + {4'b0000, e2[108]}%3329;
                                                                                                                                                                                     result[1][109] = decom_out[1][109]+ mul_add_t[1][109] + {4'b0000, e2[109]}%3329;
                                                                                                                                                                                     result[1][110] = decom_out[1][110]+ mul_add_t[1][110] + {4'b0000, e2[110]}%3329;
                                                                                                                                                                                     result[1][111] = decom_out[1][111]+ mul_add_t[1][111] + {4'b0000, e2[111]}%3329;
                                                                                                                                                                                     result[1][112] = decom_out[1][112]+ mul_add_t[1][112] + {4'b0000, e2[112]}%3329;
                                                                                                                                                                                     result[1][113] = decom_out[1][113]+ mul_add_t[1][113] + {4'b0000, e2[113]}%3329;
                                                                                                                                                                                     result[1][114] = decom_out[1][114]+ mul_add_t[1][114] + {4'b0000, e2[114]}%3329;
                                                                                                                                                                                     result[1][115] = decom_out[1][115]+ mul_add_t[1][115] + {4'b0000, e2[115]}%3329;
                                                                                                                                                                                     result[1][116] = decom_out[1][116]+ mul_add_t[1][116] + {4'b0000, e2[116]}%3329;
                                                                                                                                                                                     result[1][117] = decom_out[1][117]+ mul_add_t[1][117] + {4'b0000, e2[117]}%3329;
                                                                                                                                                                                     result[1][118] = decom_out[1][118]+ mul_add_t[1][118] + {4'b0000, e2[118]}%3329;
                                                                                                                                                                                     result[1][119] = decom_out[1][119]+ mul_add_t[1][119] + {4'b0000, e2[119]}%3329;
                                                                                                                                                                                     result[1][120] = decom_out[1][120]+ mul_add_t[1][120] + {4'b0000, e2[120]}%3329;
                                                                                                                                                                                     result[1][121] = decom_out[1][121]+ mul_add_t[1][121] + {4'b0000, e2[121]}%3329;
                                                                                                                                                                                     result[1][122] = decom_out[1][122]+ mul_add_t[1][122] + {4'b0000, e2[122]}%3329;
                                                                                                                                                                                     result[1][123] = decom_out[1][123]+ mul_add_t[1][123] + {4'b0000, e2[123]}%3329;
                                                                                                                                                                                     result[1][124] = decom_out[1][124]+ mul_add_t[1][124] + {4'b0000, e2[124]}%3329;
                                                                                                                                                                                     result[1][125] = decom_out[1][125]+ mul_add_t[1][125] + {4'b0000, e2[125]}%3329;
                                                                                                                                                                                     result[1][126] = decom_out[1][126]+ mul_add_t[1][126] + {4'b0000, e2[126]}%3329;
                                                                                                                                                                                     result[1][127] = decom_out[1][127]+ mul_add_t[1][127] + {4'b0000, e2[127]}%3329;
                                                                                                                                                                                     result[1][128] = decom_out[1][128]+ mul_add_t[1][128] + {4'b0000, e2[128]}%3329;
                                                                                                                                                                                     result[1][129] = decom_out[1][129]+ mul_add_t[1][129] + {4'b0000, e2[129]}%3329;
                                                                                                                                                                                     result[1][130] = decom_out[1][130]+ mul_add_t[1][130] + {4'b0000, e2[130]}%3329;
                                                                                                                                                                                     result[1][131] = decom_out[1][131]+ mul_add_t[1][131] + {4'b0000, e2[131]}%3329;
                                                                                                                                                                                     result[1][132] = decom_out[1][132]+ mul_add_t[1][132] + {4'b0000, e2[132]}%3329;
                                                                                                                                                                                     result[1][133] = decom_out[1][133]+ mul_add_t[1][133] + {4'b0000, e2[133]}%3329;
                                                                                                                                                                                     result[1][134] = decom_out[1][134]+ mul_add_t[1][134] + {4'b0000, e2[134]}%3329;
                                                                                                                                                                                     result[1][135] = decom_out[1][135]+ mul_add_t[1][135] + {4'b0000, e2[135]}%3329;
                                                                                                                                                                                     result[1][136] = decom_out[1][136]+ mul_add_t[1][136] + {4'b0000, e2[136]}%3329;
                                                                                                                                                                                     result[1][137] = decom_out[1][137]+ mul_add_t[1][137] + {4'b0000, e2[137]}%3329;
                                                                                                                                                                                     result[1][138] = decom_out[1][138]+ mul_add_t[1][138] + {4'b0000, e2[138]}%3329;
                                                                                                                                                                                     result[1][139] = decom_out[1][139]+ mul_add_t[1][139] + {4'b0000, e2[139]}%3329;
                                                                                                                                                                                     result[1][140] = decom_out[1][140]+ mul_add_t[1][140] + {4'b0000, e2[140]}%3329;
                                                                                                                                                                                     result[1][141] = decom_out[1][141]+ mul_add_t[1][141] + {4'b0000, e2[141]}%3329;
                                                                                                                                                                                     result[1][142] = decom_out[1][142]+ mul_add_t[1][142] + {4'b0000, e2[142]}%3329;
                                                                                                                                                                                     result[1][143] = decom_out[1][143]+ mul_add_t[1][143] + {4'b0000, e2[143]}%3329;
                                                                                                                                                                                     result[1][144] = decom_out[1][144]+ mul_add_t[1][144] + {4'b0000, e2[144]}%3329;
                                                                                                                                                                                     result[1][145] = decom_out[1][145]+ mul_add_t[1][145] + {4'b0000, e2[145]}%3329;
                                                                                                                                                                                     result[1][146] = decom_out[1][146]+ mul_add_t[1][146] + {4'b0000, e2[146]}%3329;
                                                                                                                                                                                     result[1][147] = decom_out[1][147]+ mul_add_t[1][147] + {4'b0000, e2[147]}%3329;
                                                                                                                                                                                     result[1][148] = decom_out[1][148]+ mul_add_t[1][148] + {4'b0000, e2[148]}%3329;
                                                                                                                                                                                     result[1][149] = decom_out[1][149]+ mul_add_t[1][149] + {4'b0000, e2[149]}%3329;
                                                                                                                                                                                     result[1][150] = decom_out[1][150]+ mul_add_t[1][150] + {4'b0000, e2[150]}%3329;
                                                                                                                                                                                     result[1][151] = decom_out[1][151]+ mul_add_t[1][151] + {4'b0000, e2[151]}%3329;
                                                                                                                                                                                     result[1][152] = decom_out[1][152]+ mul_add_t[1][152] + {4'b0000, e2[152]}%3329;
                                                                                                                                                                                     result[1][153] = decom_out[1][153]+ mul_add_t[1][153] + {4'b0000, e2[153]}%3329;
                                                                                                                                                                                     result[1][154] = decom_out[1][154]+ mul_add_t[1][154] + {4'b0000, e2[154]}%3329;
                                                                                                                                                                                     result[1][155] = decom_out[1][155]+ mul_add_t[1][155] + {4'b0000, e2[155]}%3329;
                                                                                                                                                                                     result[1][156] = decom_out[1][156]+ mul_add_t[1][156] + {4'b0000, e2[156]}%3329;
                                                                                                                                                                                     result[1][157] = decom_out[1][157]+ mul_add_t[1][157] + {4'b0000, e2[157]}%3329;
                                                                                                                                                                                     result[1][158] = decom_out[1][158]+ mul_add_t[1][158] + {4'b0000, e2[158]}%3329;
                                                                                                                                                                                     result[1][159] = decom_out[1][159]+ mul_add_t[1][159] + {4'b0000, e2[159]}%3329;
                                                                                                                                                                                     result[1][160] = decom_out[1][160]+ mul_add_t[1][160] + {4'b0000, e2[160]}%3329;
                                                                                                                                                                                     result[1][161] = decom_out[1][161]+ mul_add_t[1][161] + {4'b0000, e2[161]}%3329;
                                                                                                                                                                                     result[1][162] = decom_out[1][162]+ mul_add_t[1][162] + {4'b0000, e2[162]}%3329;
                                                                                                                                                                                     result[1][163] = decom_out[1][163]+ mul_add_t[1][163] + {4'b0000, e2[163]}%3329;
                                                                                                                                                                                     result[1][164] = decom_out[1][164]+ mul_add_t[1][164] + {4'b0000, e2[164]}%3329;
                                                                                                                                                                                     result[1][165] = decom_out[1][165]+ mul_add_t[1][165] + {4'b0000, e2[165]}%3329;
                                                                                                                                                                                     result[1][166] = decom_out[1][166]+ mul_add_t[1][166] + {4'b0000, e2[166]}%3329;
                                                                                                                                                                                     result[1][167] = decom_out[1][167]+ mul_add_t[1][167] + {4'b0000, e2[167]}%3329;
                                                                                                                                                                                     result[1][168] = decom_out[1][168]+ mul_add_t[1][168] + {4'b0000, e2[168]}%3329;
                                                                                                                                                                                     result[1][169] = decom_out[1][169]+ mul_add_t[1][169] + {4'b0000, e2[169]}%3329;
                                                                                                                                                                                     result[1][170] = decom_out[1][170]+ mul_add_t[1][170] + {4'b0000, e2[170]}%3329;
                                                                                                                                                                                     result[1][171] = decom_out[1][171]+ mul_add_t[1][171] + {4'b0000, e2[171]}%3329;
                                                                                                                                                                                     result[1][172] = decom_out[1][172]+ mul_add_t[1][172] + {4'b0000, e2[172]}%3329;
                                                                                                                                                                                     result[1][173] = decom_out[1][173]+ mul_add_t[1][173] + {4'b0000, e2[173]}%3329;
                                                                                                                                                                                     result[1][174] = decom_out[1][174]+ mul_add_t[1][174] + {4'b0000, e2[174]}%3329;
                                                                                                                                                                                     result[1][175] = decom_out[1][175]+ mul_add_t[1][175] + {4'b0000, e2[175]}%3329;
                                                                                                                                                                                     result[1][176] = decom_out[1][176]+ mul_add_t[1][176] + {4'b0000, e2[176]}%3329;
                                                                                                                                                                                     result[1][177] = decom_out[1][177]+ mul_add_t[1][177] + {4'b0000, e2[177]}%3329;
                                                                                                                                                                                     result[1][178] = decom_out[1][178]+ mul_add_t[1][178] + {4'b0000, e2[178]}%3329;
                                                                                                                                                                                     result[1][179] = decom_out[1][179]+ mul_add_t[1][179] + {4'b0000, e2[179]}%3329;
                                                                                                                                                                                     result[1][180] = decom_out[1][180]+ mul_add_t[1][180] + {4'b0000, e2[180]}%3329;
                                                                                                                                                                                     result[1][181] = decom_out[1][181]+ mul_add_t[1][181] + {4'b0000, e2[181]}%3329;
                                                                                                                                                                                     result[1][182] = decom_out[1][182]+ mul_add_t[1][182] + {4'b0000, e2[182]}%3329;
                                                                                                                                                                                     result[1][183] = decom_out[1][183]+ mul_add_t[1][183] + {4'b0000, e2[183]}%3329;
                                                                                                                                                                                     result[1][184] = decom_out[1][184]+ mul_add_t[1][184] + {4'b0000, e2[184]}%3329;
                                                                                                                                                                                     result[1][185] = decom_out[1][185]+ mul_add_t[1][185] + {4'b0000, e2[185]}%3329;
                                                                                                                                                                                     result[1][186] = decom_out[1][186]+ mul_add_t[1][186] + {4'b0000, e2[186]}%3329;
                                                                                                                                                                                     result[1][187] = decom_out[1][187]+ mul_add_t[1][187] + {4'b0000, e2[187]}%3329;
                                                                                                                                                                                     result[1][188] = decom_out[1][188]+ mul_add_t[1][188] + {4'b0000, e2[188]}%3329;
                                                                                                                                                                                     result[1][189] = decom_out[1][189]+ mul_add_t[1][189] + {4'b0000, e2[189]}%3329;
                                                                                                                                                                                     result[1][190] = decom_out[1][190]+ mul_add_t[1][190] + {4'b0000, e2[190]}%3329;
                                                                                                                                                                                     result[1][191] = decom_out[1][191]+ mul_add_t[1][191] + {4'b0000, e2[191]}%3329;
                                                                                                                                                                                     result[1][192] = decom_out[1][192]+ mul_add_t[1][192] + {4'b0000, e2[192]}%3329;
                                                                                                                                                                                     result[1][193] = decom_out[1][193]+ mul_add_t[1][193] + {4'b0000, e2[193]}%3329;
                                                                                                                                                                                     result[1][194] = decom_out[1][194]+ mul_add_t[1][194] + {4'b0000, e2[194]}%3329;
                                                                                                                                                                                     result[1][195] = decom_out[1][195]+ mul_add_t[1][195] + {4'b0000, e2[195]}%3329;
                                                                                                                                                                                     result[1][196] = decom_out[1][196]+ mul_add_t[1][196] + {4'b0000, e2[196]}%3329;
                                                                                                                                                                                     result[1][197] = decom_out[1][197]+ mul_add_t[1][197] + {4'b0000, e2[197]}%3329;
                                                                                                                                                                                     result[1][198] = decom_out[1][198]+ mul_add_t[1][198] + {4'b0000, e2[198]}%3329;
                                                                                                                                                                                     result[1][199] = decom_out[1][199]+ mul_add_t[1][199] + {4'b0000, e2[199]}%3329;
                                                                                                                                                                                     result[1][200] = decom_out[1][200]+ mul_add_t[1][200] + {4'b0000, e2[200]}%3329;
                                                                                                                                                                                     result[1][201] = decom_out[1][201]+ mul_add_t[1][201] + {4'b0000, e2[201]}%3329;
                                                                                                                                                                                     result[1][202] = decom_out[1][202]+ mul_add_t[1][202] + {4'b0000, e2[202]}%3329;
                                                                                                                                                                                     result[1][203] = decom_out[1][203]+ mul_add_t[1][203] + {4'b0000, e2[203]}%3329;
                                                                                                                                                                                     result[1][204] = decom_out[1][204]+ mul_add_t[1][204] + {4'b0000, e2[204]}%3329;
                                                                                                                                                                                     result[1][205] = decom_out[1][205]+ mul_add_t[1][205] + {4'b0000, e2[205]}%3329;
                                                                                                                                                                                     result[1][206] = decom_out[1][206]+ mul_add_t[1][206] + {4'b0000, e2[206]}%3329;
                                                                                                                                                                                     result[1][207] = decom_out[1][207]+ mul_add_t[1][207] + {4'b0000, e2[207]}%3329;
                                                                                                                                                                                     result[1][208] = decom_out[1][208]+ mul_add_t[1][208] + {4'b0000, e2[208]}%3329;
                                                                                                                                                                                     result[1][209] = decom_out[1][209]+ mul_add_t[1][209] + {4'b0000, e2[209]}%3329;
                                                                                                                                                                                     result[1][210] = decom_out[1][210]+ mul_add_t[1][210] + {4'b0000, e2[210]}%3329;
                                                                                                                                                                                     result[1][211] = decom_out[1][211]+ mul_add_t[1][211] + {4'b0000, e2[211]}%3329;
                                                                                                                                                                                     result[1][212] = decom_out[1][212]+ mul_add_t[1][212] + {4'b0000, e2[212]}%3329;
                                                                                                                                                                                     result[1][213] = decom_out[1][213]+ mul_add_t[1][213] + {4'b0000, e2[213]}%3329;
                                                                                                                                                                                     result[1][214] = decom_out[1][214]+ mul_add_t[1][214] + {4'b0000, e2[214]}%3329;
                                                                                                                                                                                     result[1][215] = decom_out[1][215]+ mul_add_t[1][215] + {4'b0000, e2[215]}%3329;
                                                                                                                                                                                     result[1][216] = decom_out[1][216]+ mul_add_t[1][216] + {4'b0000, e2[216]}%3329;
                                                                                                                                                                                     result[1][217] = decom_out[1][217]+ mul_add_t[1][217] + {4'b0000, e2[217]}%3329;
                                                                                                                                                                                     result[1][218] = decom_out[1][218]+ mul_add_t[1][218] + {4'b0000, e2[218]}%3329;
                                                                                                                                                                                     result[1][219] = decom_out[1][219]+ mul_add_t[1][219] + {4'b0000, e2[219]}%3329;
                                                                                                                                                                                     result[1][220] = decom_out[1][220]+ mul_add_t[1][220] + {4'b0000, e2[220]}%3329;
                                                                                                                                                                                     result[1][221] = decom_out[1][221]+ mul_add_t[1][221] + {4'b0000, e2[221]}%3329;
                                                                                                                                                                                     result[1][222] = decom_out[1][222]+ mul_add_t[1][222] + {4'b0000, e2[222]}%3329;
                                                                                                                                                                                     result[1][223] = decom_out[1][223]+ mul_add_t[1][223] + {4'b0000, e2[223]}%3329;
                                                                                                                                                                                     result[1][224] = decom_out[1][224]+ mul_add_t[1][224] + {4'b0000, e2[224]}%3329;
                                                                                                                                                                                     result[1][225] = decom_out[1][225]+ mul_add_t[1][225] + {4'b0000, e2[225]}%3329;
                                                                                                                                                                                     result[1][226] = decom_out[1][226]+ mul_add_t[1][226] + {4'b0000, e2[226]}%3329;
                                                                                                                                                                                     result[1][227] = decom_out[1][227]+ mul_add_t[1][227] + {4'b0000, e2[227]}%3329;
                                                                                                                                                                                     result[1][228] = decom_out[1][228]+ mul_add_t[1][228] + {4'b0000, e2[228]}%3329;
                                                                                                                                                                                     result[1][229] = decom_out[1][229]+ mul_add_t[1][229] + {4'b0000, e2[229]}%3329;
                                                                                                                                                                                     result[1][230] = decom_out[1][230]+ mul_add_t[1][230] + {4'b0000, e2[230]}%3329;
                                                                                                                                                                                     result[1][231] = decom_out[1][231]+ mul_add_t[1][231] + {4'b0000, e2[231]}%3329;
                                                                                                                                                                                     result[1][232] = decom_out[1][232]+ mul_add_t[1][232] + {4'b0000, e2[232]}%3329;
                                                                                                                                                                                     result[1][233] = decom_out[1][233]+ mul_add_t[1][233] + {4'b0000, e2[233]}%3329;
                                                                                                                                                                                     result[1][234] = decom_out[1][234]+ mul_add_t[1][234] + {4'b0000, e2[234]}%3329;
                                                                                                                                                                                     result[1][235] = decom_out[1][235]+ mul_add_t[1][235] + {4'b0000, e2[235]}%3329;
                                                                                                                                                                                     result[1][236] = decom_out[1][236]+ mul_add_t[1][236] + {4'b0000, e2[236]}%3329;
                                                                                                                                                                                     result[1][237] = decom_out[1][237]+ mul_add_t[1][237] + {4'b0000, e2[237]}%3329;
                                                                                                                                                                                     result[1][238] = decom_out[1][238]+ mul_add_t[1][238] + {4'b0000, e2[238]}%3329;
                                                                                                                                                                                     result[1][239] = decom_out[1][239]+ mul_add_t[1][239] + {4'b0000, e2[239]}%3329;
                                                                                                                                                                                     result[1][240] = decom_out[1][240]+ mul_add_t[1][240] + {4'b0000, e2[240]}%3329;
                                                                                                                                                                                     result[1][241] = decom_out[1][241]+ mul_add_t[1][241] + {4'b0000, e2[241]}%3329;
                                                                                                                                                                                     result[1][242] = decom_out[1][242]+ mul_add_t[1][242] + {4'b0000, e2[242]}%3329;
                                                                                                                                                                                     result[1][243] = decom_out[1][243]+ mul_add_t[1][243] + {4'b0000, e2[243]}%3329;
                                                                                                                                                                                     result[1][244] = decom_out[1][244]+ mul_add_t[1][244] + {4'b0000, e2[244]}%3329;
                                                                                                                                                                                     result[1][245] = decom_out[1][245]+ mul_add_t[1][245] + {4'b0000, e2[245]}%3329;
                                                                                                                                                                                     result[1][246] = decom_out[1][246]+ mul_add_t[1][246] + {4'b0000, e2[246]}%3329;
                                                                                                                                                                                     result[1][247] = decom_out[1][247]+ mul_add_t[1][247] + {4'b0000, e2[247]}%3329;
                                                                                                                                                                                     result[1][248] = decom_out[1][248]+ mul_add_t[1][248] + {4'b0000, e2[248]}%3329;
                                                                                                                                                                                     result[1][249] = decom_out[1][249]+ mul_add_t[1][249] + {4'b0000, e2[249]}%3329;
                                                                                                                                                                                     result[1][250] = decom_out[1][250]+ mul_add_t[1][250] + {4'b0000, e2[250]}%3329;
                                                                                                                                                                                     result[1][251] = decom_out[1][251]+ mul_add_t[1][251] + {4'b0000, e2[251]}%3329;
                                                                                                                                                                                     result[1][252] = decom_out[1][252]+ mul_add_t[1][252] + {4'b0000, e2[252]}%3329;
                                                                                                                                                                                     result[1][253] = decom_out[1][253]+ mul_add_t[1][253] + {4'b0000, e2[253]}%3329;
                                                                                                                                                                                     result[1][254] = decom_out[1][254]+ mul_add_t[1][254] + {4'b0000, e2[254]}%3329;
                                                                                                                                                                                     result[1][255] = decom_out[1][255]+ mul_add_t[1][255] + {4'b0000, e2[255]}%3329;
                                                                                                                                                                                     result[2][0] = decom_out[2][0]+ mul_add_t[2][0] + {4'b0000, e2[0]}%3329;
                                                                                                                                                                                     result[2][1] = decom_out[2][1]+ mul_add_t[2][1] + {4'b0000, e2[1]}%3329;
                                                                                                                                                                                     result[2][2] = decom_out[2][2]+ mul_add_t[2][2] + {4'b0000, e2[2]}%3329;
                                                                                                                                                                                     result[2][3] = decom_out[2][3]+ mul_add_t[2][3] + {4'b0000, e2[3]}%3329;
                                                                                                                                                                                     result[2][4] = decom_out[2][4]+ mul_add_t[2][4] + {4'b0000, e2[4]}%3329;
                                                                                                                                                                                     result[2][5] = decom_out[2][5]+ mul_add_t[2][5] + {4'b0000, e2[5]}%3329;
                                                                                                                                                                                     result[2][6] = decom_out[2][6]+ mul_add_t[2][6] + {4'b0000, e2[6]}%3329;
                                                                                                                                                                                     result[2][7] = decom_out[2][7]+ mul_add_t[2][7] + {4'b0000, e2[7]}%3329;
                                                                                                                                                                                     result[2][8] = decom_out[2][8]+ mul_add_t[2][8] + {4'b0000, e2[8]}%3329;
                                                                                                                                                                                     result[2][9] = decom_out[2][9]+ mul_add_t[2][9] + {4'b0000, e2[9]}%3329;
                                                                                                                                                                                     result[2][10] = decom_out[2][10]+ mul_add_t[2][10] + {4'b0000, e2[10]}%3329;
                                                                                                                                                                                     result[2][11] = decom_out[2][11]+ mul_add_t[2][11] + {4'b0000, e2[11]}%3329;
                                                                                                                                                                                     result[2][12] = decom_out[2][12]+ mul_add_t[2][12] + {4'b0000, e2[12]}%3329;
                                                                                                                                                                                     result[2][13] = decom_out[2][13]+ mul_add_t[2][13] + {4'b0000, e2[13]}%3329;
                                                                                                                                                                                     result[2][14] = decom_out[2][14]+ mul_add_t[2][14] + {4'b0000, e2[14]}%3329;
                                                                                                                                                                                     result[2][15] = decom_out[2][15]+ mul_add_t[2][15] + {4'b0000, e2[15]}%3329;
                                                                                                                                                                                     result[2][16] = decom_out[2][16]+ mul_add_t[2][16] + {4'b0000, e2[16]}%3329;
                                                                                                                                                                                     result[2][17] = decom_out[2][17]+ mul_add_t[2][17] + {4'b0000, e2[17]}%3329;
                                                                                                                                                                                     result[2][18] = decom_out[2][18]+ mul_add_t[2][18] + {4'b0000, e2[18]}%3329;
                                                                                                                                                                                     result[2][19] = decom_out[2][19]+ mul_add_t[2][19] + {4'b0000, e2[19]}%3329;
                                                                                                                                                                                     result[2][20] = decom_out[2][20]+ mul_add_t[2][20] + {4'b0000, e2[20]}%3329;
                                                                                                                                                                                     result[2][21] = decom_out[2][21]+ mul_add_t[2][21] + {4'b0000, e2[21]}%3329;
                                                                                                                                                                                     result[2][22] = decom_out[2][22]+ mul_add_t[2][22] + {4'b0000, e2[22]}%3329;
                                                                                                                                                                                     result[2][23] = decom_out[2][23]+ mul_add_t[2][23] + {4'b0000, e2[23]}%3329;
                                                                                                                                                                                     result[2][24] = decom_out[2][24]+ mul_add_t[2][24] + {4'b0000, e2[24]}%3329;
                                                                                                                                                                                     result[2][25] = decom_out[2][25]+ mul_add_t[2][25] + {4'b0000, e2[25]}%3329;
                                                                                                                                                                                     result[2][26] = decom_out[2][26]+ mul_add_t[2][26] + {4'b0000, e2[26]}%3329;
                                                                                                                                                                                     result[2][27] = decom_out[2][27]+ mul_add_t[2][27] + {4'b0000, e2[27]}%3329;
                                                                                                                                                                                     result[2][28] = decom_out[2][28]+ mul_add_t[2][28] + {4'b0000, e2[28]}%3329;
                                                                                                                                                                                     result[2][29] = decom_out[2][29]+ mul_add_t[2][29] + {4'b0000, e2[29]}%3329;
                                                                                                                                                                                     result[2][30] = decom_out[2][30]+ mul_add_t[2][30] + {4'b0000, e2[30]}%3329;
                                                                                                                                                                                     result[2][31] = decom_out[2][31]+ mul_add_t[2][31] + {4'b0000, e2[31]}%3329;
                                                                                                                                                                                     result[2][32] = decom_out[2][32]+ mul_add_t[2][32] + {4'b0000, e2[32]}%3329;
                                                                                                                                                                                     result[2][33] = decom_out[2][33]+ mul_add_t[2][33] + {4'b0000, e2[33]}%3329;
                                                                                                                                                                                     result[2][34] = decom_out[2][34]+ mul_add_t[2][34] + {4'b0000, e2[34]}%3329;
                                                                                                                                                                                     result[2][35] = decom_out[2][35]+ mul_add_t[2][35] + {4'b0000, e2[35]}%3329;
                                                                                                                                                                                     result[2][36] = decom_out[2][36]+ mul_add_t[2][36] + {4'b0000, e2[36]}%3329;
                                                                                                                                                                                     result[2][37] = decom_out[2][37]+ mul_add_t[2][37] + {4'b0000, e2[37]}%3329;
                                                                                                                                                                                     result[2][38] = decom_out[2][38]+ mul_add_t[2][38] + {4'b0000, e2[38]}%3329;
                                                                                                                                                                                     result[2][39] = decom_out[2][39]+ mul_add_t[2][39] + {4'b0000, e2[39]}%3329;
                                                                                                                                                                                     result[2][40] = decom_out[2][40]+ mul_add_t[2][40] + {4'b0000, e2[40]}%3329;
                                                                                                                                                                                     result[2][41] = decom_out[2][41]+ mul_add_t[2][41] + {4'b0000, e2[41]}%3329;
                                                                                                                                                                                     result[2][42] = decom_out[2][42]+ mul_add_t[2][42] + {4'b0000, e2[42]}%3329;
                                                                                                                                                                                     result[2][43] = decom_out[2][43]+ mul_add_t[2][43] + {4'b0000, e2[43]}%3329;
                                                                                                                                                                                     result[2][44] = decom_out[2][44]+ mul_add_t[2][44] + {4'b0000, e2[44]}%3329;
                                                                                                                                                                                     result[2][45] = decom_out[2][45]+ mul_add_t[2][45] + {4'b0000, e2[45]}%3329;
                                                                                                                                                                                     result[2][46] = decom_out[2][46]+ mul_add_t[2][46] + {4'b0000, e2[46]}%3329;
                                                                                                                                                                                     result[2][47] = decom_out[2][47]+ mul_add_t[2][47] + {4'b0000, e2[47]}%3329;
                                                                                                                                                                                     result[2][48] = decom_out[2][48]+ mul_add_t[2][48] + {4'b0000, e2[48]}%3329;
                                                                                                                                                                                     result[2][49] = decom_out[2][49]+ mul_add_t[2][49] + {4'b0000, e2[49]}%3329;
                                                                                                                                                                                     result[2][50] = decom_out[2][50]+ mul_add_t[2][50] + {4'b0000, e2[50]}%3329;
                                                                                                                                                                                     result[2][51] = decom_out[2][51]+ mul_add_t[2][51] + {4'b0000, e2[51]}%3329;
                                                                                                                                                                                     result[2][52] = decom_out[2][52]+ mul_add_t[2][52] + {4'b0000, e2[52]}%3329;
                                                                                                                                                                                     result[2][53] = decom_out[2][53]+ mul_add_t[2][53] + {4'b0000, e2[53]}%3329;
                                                                                                                                                                                     result[2][54] = decom_out[2][54]+ mul_add_t[2][54] + {4'b0000, e2[54]}%3329;
                                                                                                                                                                                     result[2][55] = decom_out[2][55]+ mul_add_t[2][55] + {4'b0000, e2[55]}%3329;
                                                                                                                                                                                     result[2][56] = decom_out[2][56]+ mul_add_t[2][56] + {4'b0000, e2[56]}%3329;
                                                                                                                                                                                     result[2][57] = decom_out[2][57]+ mul_add_t[2][57] + {4'b0000, e2[57]}%3329;
                                                                                                                                                                                     result[2][58] = decom_out[2][58]+ mul_add_t[2][58] + {4'b0000, e2[58]}%3329;
                                                                                                                                                                                     result[2][59] = decom_out[2][59]+ mul_add_t[2][59] + {4'b0000, e2[59]}%3329;
                                                                                                                                                                                     result[2][60] = decom_out[2][60]+ mul_add_t[2][60] + {4'b0000, e2[60]}%3329;
                                                                                                                                                                                     result[2][61] = decom_out[2][61]+ mul_add_t[2][61] + {4'b0000, e2[61]}%3329;
                                                                                                                                                                                     result[2][62] = decom_out[2][62]+ mul_add_t[2][62] + {4'b0000, e2[62]}%3329;
                                                                                                                                                                                     result[2][63] = decom_out[2][63]+ mul_add_t[2][63] + {4'b0000, e2[63]}%3329;
                                                                                                                                                                                     result[2][64] = decom_out[2][64]+ mul_add_t[2][64] + {4'b0000, e2[64]}%3329;
                                                                                                                                                                                     result[2][65] = decom_out[2][65]+ mul_add_t[2][65] + {4'b0000, e2[65]}%3329;
                                                                                                                                                                                     result[2][66] = decom_out[2][66]+ mul_add_t[2][66] + {4'b0000, e2[66]}%3329;
                                                                                                                                                                                     result[2][67] = decom_out[2][67]+ mul_add_t[2][67] + {4'b0000, e2[67]}%3329;
                                                                                                                                                                                     result[2][68] = decom_out[2][68]+ mul_add_t[2][68] + {4'b0000, e2[68]}%3329;
                                                                                                                                                                                     result[2][69] = decom_out[2][69]+ mul_add_t[2][69] + {4'b0000, e2[69]}%3329;
                                                                                                                                                                                     result[2][70] = decom_out[2][70]+ mul_add_t[2][70] + {4'b0000, e2[70]}%3329;
                                                                                                                                                                                     result[2][71] = decom_out[2][71]+ mul_add_t[2][71] + {4'b0000, e2[71]}%3329;
                                                                                                                                                                                     result[2][72] = decom_out[2][72]+ mul_add_t[2][72] + {4'b0000, e2[72]}%3329;
                                                                                                                                                                                     result[2][73] = decom_out[2][73]+ mul_add_t[2][73] + {4'b0000, e2[73]}%3329;
                                                                                                                                                                                     result[2][74] = decom_out[2][74]+ mul_add_t[2][74] + {4'b0000, e2[74]}%3329;
                                                                                                                                                                                     result[2][75] = decom_out[2][75]+ mul_add_t[2][75] + {4'b0000, e2[75]}%3329;
                                                                                                                                                                                     result[2][76] = decom_out[2][76]+ mul_add_t[2][76] + {4'b0000, e2[76]}%3329;
                                                                                                                                                                                     result[2][77] = decom_out[2][77]+ mul_add_t[2][77] + {4'b0000, e2[77]}%3329;
                                                                                                                                                                                     result[2][78] = decom_out[2][78]+ mul_add_t[2][78] + {4'b0000, e2[78]}%3329;
                                                                                                                                                                                     result[2][79] = decom_out[2][79]+ mul_add_t[2][79] + {4'b0000, e2[79]}%3329;
                                                                                                                                                                                     result[2][80] = decom_out[2][80]+ mul_add_t[2][80] + {4'b0000, e2[80]}%3329;
                                                                                                                                                                                     result[2][81] = decom_out[2][81]+ mul_add_t[2][81] + {4'b0000, e2[81]}%3329;
                                                                                                                                                                                     result[2][82] = decom_out[2][82]+ mul_add_t[2][82] + {4'b0000, e2[82]}%3329;
                                                                                                                                                                                     result[2][83] = decom_out[2][83]+ mul_add_t[2][83] + {4'b0000, e2[83]}%3329;
                                                                                                                                                                                     result[2][84] = decom_out[2][84]+ mul_add_t[2][84] + {4'b0000, e2[84]}%3329;
                                                                                                                                                                                     result[2][85] = decom_out[2][85]+ mul_add_t[2][85] + {4'b0000, e2[85]}%3329;
                                                                                                                                                                                     result[2][86] = decom_out[2][86]+ mul_add_t[2][86] + {4'b0000, e2[86]}%3329;
                                                                                                                                                                                     result[2][87] = decom_out[2][87]+ mul_add_t[2][87] + {4'b0000, e2[87]}%3329;
                                                                                                                                                                                     result[2][88] = decom_out[2][88]+ mul_add_t[2][88] + {4'b0000, e2[88]}%3329;
                                                                                                                                                                                     result[2][89] = decom_out[2][89]+ mul_add_t[2][89] + {4'b0000, e2[89]}%3329;
                                                                                                                                                                                     result[2][90] = decom_out[2][90]+ mul_add_t[2][90] + {4'b0000, e2[90]}%3329;
                                                                                                                                                                                     result[2][91] = decom_out[2][91]+ mul_add_t[2][91] + {4'b0000, e2[91]}%3329;
                                                                                                                                                                                     result[2][92] = decom_out[2][92]+ mul_add_t[2][92] + {4'b0000, e2[92]}%3329;
                                                                                                                                                                                     result[2][93] = decom_out[2][93]+ mul_add_t[2][93] + {4'b0000, e2[93]}%3329;
                                                                                                                                                                                     result[2][94] = decom_out[2][94]+ mul_add_t[2][94] + {4'b0000, e2[94]}%3329;
                                                                                                                                                                                     result[2][95] = decom_out[2][95]+ mul_add_t[2][95] + {4'b0000, e2[95]}%3329;
                                                                                                                                                                                     result[2][96] = decom_out[2][96]+ mul_add_t[2][96] + {4'b0000, e2[96]}%3329;
                                                                                                                                                                                     result[2][97] = decom_out[2][97]+ mul_add_t[2][97] + {4'b0000, e2[97]}%3329;
                                                                                                                                                                                     result[2][98] = decom_out[2][98]+ mul_add_t[2][98] + {4'b0000, e2[98]}%3329;
                                                                                                                                                                                     result[2][99] = decom_out[2][99]+ mul_add_t[2][99] + {4'b0000, e2[99]}%3329;
                                                                                                                                                                                     result[2][100] = decom_out[2][100]+ mul_add_t[2][100] + {4'b0000, e2[100]}%3329;
                                                                                                                                                                                     result[2][101] = decom_out[2][101]+ mul_add_t[2][101] + {4'b0000, e2[101]}%3329;
                                                                                                                                                                                     result[2][102] = decom_out[2][102]+ mul_add_t[2][102] + {4'b0000, e2[102]}%3329;
                                                                                                                                                                                     result[2][103] = decom_out[2][103]+ mul_add_t[2][103] + {4'b0000, e2[103]}%3329;
                                                                                                                                                                                     result[2][104] = decom_out[2][104]+ mul_add_t[2][104] + {4'b0000, e2[104]}%3329;
                                                                                                                                                                                     result[2][105] = decom_out[2][105]+ mul_add_t[2][105] + {4'b0000, e2[105]}%3329;
                                                                                                                                                                                     result[2][106] = decom_out[2][106]+ mul_add_t[2][106] + {4'b0000, e2[106]}%3329;
                                                                                                                                                                                     result[2][107] = decom_out[2][107]+ mul_add_t[2][107] + {4'b0000, e2[107]}%3329;
                                                                                                                                                                                     result[2][108] = decom_out[2][108]+ mul_add_t[2][108] + {4'b0000, e2[108]}%3329;
                                                                                                                                                                                     result[2][109] = decom_out[2][109]+ mul_add_t[2][109] + {4'b0000, e2[109]}%3329;
                                                                                                                                                                                     result[2][110] = decom_out[2][110]+ mul_add_t[2][110] + {4'b0000, e2[110]}%3329;
                                                                                                                                                                                     result[2][111] = decom_out[2][111]+ mul_add_t[2][111] + {4'b0000, e2[111]}%3329;
                                                                                                                                                                                     result[2][112] = decom_out[2][112]+ mul_add_t[2][112] + {4'b0000, e2[112]}%3329;
                                                                                                                                                                                     result[2][113] = decom_out[2][113]+ mul_add_t[2][113] + {4'b0000, e2[113]}%3329;
                                                                                                                                                                                     result[2][114] = decom_out[2][114]+ mul_add_t[2][114] + {4'b0000, e2[114]}%3329;
                                                                                                                                                                                     result[2][115] = decom_out[2][115]+ mul_add_t[2][115] + {4'b0000, e2[115]}%3329;
                                                                                                                                                                                     result[2][116] = decom_out[2][116]+ mul_add_t[2][116] + {4'b0000, e2[116]}%3329;
                                                                                                                                                                                     result[2][117] = decom_out[2][117]+ mul_add_t[2][117] + {4'b0000, e2[117]}%3329;
                                                                                                                                                                                     result[2][118] = decom_out[2][118]+ mul_add_t[2][118] + {4'b0000, e2[118]}%3329;
                                                                                                                                                                                     result[2][119] = decom_out[2][119]+ mul_add_t[2][119] + {4'b0000, e2[119]}%3329;
                                                                                                                                                                                     result[2][120] = decom_out[2][120]+ mul_add_t[2][120] + {4'b0000, e2[120]}%3329;
                                                                                                                                                                                     result[2][121] = decom_out[2][121]+ mul_add_t[2][121] + {4'b0000, e2[121]}%3329;
                                                                                                                                                                                     result[2][122] = decom_out[2][122]+ mul_add_t[2][122] + {4'b0000, e2[122]}%3329;
                                                                                                                                                                                     result[2][123] = decom_out[2][123]+ mul_add_t[2][123] + {4'b0000, e2[123]}%3329;
                                                                                                                                                                                     result[2][124] = decom_out[2][124]+ mul_add_t[2][124] + {4'b0000, e2[124]}%3329;
                                                                                                                                                                                     result[2][125] = decom_out[2][125]+ mul_add_t[2][125] + {4'b0000, e2[125]}%3329;
                                                                                                                                                                                     result[2][126] = decom_out[2][126]+ mul_add_t[2][126] + {4'b0000, e2[126]}%3329;
                                                                                                                                                                                     result[2][127] = decom_out[2][127]+ mul_add_t[2][127] + {4'b0000, e2[127]}%3329;
                                                                                                                                                                                     result[2][128] = decom_out[2][128]+ mul_add_t[2][128] + {4'b0000, e2[128]}%3329;
                                                                                                                                                                                     result[2][129] = decom_out[2][129]+ mul_add_t[2][129] + {4'b0000, e2[129]}%3329;
                                                                                                                                                                                     result[2][130] = decom_out[2][130]+ mul_add_t[2][130] + {4'b0000, e2[130]}%3329;
                                                                                                                                                                                     result[2][131] = decom_out[2][131]+ mul_add_t[2][131] + {4'b0000, e2[131]}%3329;
                                                                                                                                                                                     result[2][132] = decom_out[2][132]+ mul_add_t[2][132] + {4'b0000, e2[132]}%3329;
                                                                                                                                                                                     result[2][133] = decom_out[2][133]+ mul_add_t[2][133] + {4'b0000, e2[133]}%3329;
                                                                                                                                                                                     result[2][134] = decom_out[2][134]+ mul_add_t[2][134] + {4'b0000, e2[134]}%3329;
                                                                                                                                                                                     result[2][135] = decom_out[2][135]+ mul_add_t[2][135] + {4'b0000, e2[135]}%3329;
                                                                                                                                                                                     result[2][136] = decom_out[2][136]+ mul_add_t[2][136] + {4'b0000, e2[136]}%3329;
                                                                                                                                                                                     result[2][137] = decom_out[2][137]+ mul_add_t[2][137] + {4'b0000, e2[137]}%3329;
                                                                                                                                                                                     result[2][138] = decom_out[2][138]+ mul_add_t[2][138] + {4'b0000, e2[138]}%3329;
                                                                                                                                                                                     result[2][139] = decom_out[2][139]+ mul_add_t[2][139] + {4'b0000, e2[139]}%3329;
                                                                                                                                                                                     result[2][140] = decom_out[2][140]+ mul_add_t[2][140] + {4'b0000, e2[140]}%3329;
                                                                                                                                                                                     result[2][141] = decom_out[2][141]+ mul_add_t[2][141] + {4'b0000, e2[141]}%3329;
                                                                                                                                                                                     result[2][142] = decom_out[2][142]+ mul_add_t[2][142] + {4'b0000, e2[142]}%3329;
                                                                                                                                                                                     result[2][143] = decom_out[2][143]+ mul_add_t[2][143] + {4'b0000, e2[143]}%3329;
                                                                                                                                                                                     result[2][144] = decom_out[2][144]+ mul_add_t[2][144] + {4'b0000, e2[144]}%3329;
                                                                                                                                                                                     result[2][145] = decom_out[2][145]+ mul_add_t[2][145] + {4'b0000, e2[145]}%3329;
                                                                                                                                                                                     result[2][146] = decom_out[2][146]+ mul_add_t[2][146] + {4'b0000, e2[146]}%3329;
                                                                                                                                                                                     result[2][147] = decom_out[2][147]+ mul_add_t[2][147] + {4'b0000, e2[147]}%3329;
                                                                                                                                                                                     result[2][148] = decom_out[2][148]+ mul_add_t[2][148] + {4'b0000, e2[148]}%3329;
                                                                                                                                                                                     result[2][149] = decom_out[2][149]+ mul_add_t[2][149] + {4'b0000, e2[149]}%3329;
                                                                                                                                                                                     result[2][150] = decom_out[2][150]+ mul_add_t[2][150] + {4'b0000, e2[150]}%3329;
                                                                                                                                                                                     result[2][151] = decom_out[2][151]+ mul_add_t[2][151] + {4'b0000, e2[151]}%3329;
                                                                                                                                                                                     result[2][152] = decom_out[2][152]+ mul_add_t[2][152] + {4'b0000, e2[152]}%3329;
                                                                                                                                                                                     result[2][153] = decom_out[2][153]+ mul_add_t[2][153] + {4'b0000, e2[153]}%3329;
                                                                                                                                                                                     result[2][154] = decom_out[2][154]+ mul_add_t[2][154] + {4'b0000, e2[154]}%3329;
                                                                                                                                                                                     result[2][155] = decom_out[2][155]+ mul_add_t[2][155] + {4'b0000, e2[155]}%3329;
                                                                                                                                                                                     result[2][156] = decom_out[2][156]+ mul_add_t[2][156] + {4'b0000, e2[156]}%3329;
                                                                                                                                                                                     result[2][157] = decom_out[2][157]+ mul_add_t[2][157] + {4'b0000, e2[157]}%3329;
                                                                                                                                                                                     result[2][158] = decom_out[2][158]+ mul_add_t[2][158] + {4'b0000, e2[158]}%3329;
                                                                                                                                                                                     result[2][159] = decom_out[2][159]+ mul_add_t[2][159] + {4'b0000, e2[159]}%3329;
                                                                                                                                                                                     result[2][160] = decom_out[2][160]+ mul_add_t[2][160] + {4'b0000, e2[160]}%3329;
                                                                                                                                                                                     result[2][161] = decom_out[2][161]+ mul_add_t[2][161] + {4'b0000, e2[161]}%3329;
                                                                                                                                                                                     result[2][162] = decom_out[2][162]+ mul_add_t[2][162] + {4'b0000, e2[162]}%3329;
                                                                                                                                                                                     result[2][163] = decom_out[2][163]+ mul_add_t[2][163] + {4'b0000, e2[163]}%3329;
                                                                                                                                                                                     result[2][164] = decom_out[2][164]+ mul_add_t[2][164] + {4'b0000, e2[164]}%3329;
                                                                                                                                                                                     result[2][165] = decom_out[2][165]+ mul_add_t[2][165] + {4'b0000, e2[165]}%3329;
                                                                                                                                                                                     result[2][166] = decom_out[2][166]+ mul_add_t[2][166] + {4'b0000, e2[166]}%3329;
                                                                                                                                                                                     result[2][167] = decom_out[2][167]+ mul_add_t[2][167] + {4'b0000, e2[167]}%3329;
                                                                                                                                                                                     result[2][168] = decom_out[2][168]+ mul_add_t[2][168] + {4'b0000, e2[168]}%3329;
                                                                                                                                                                                     result[2][169] = decom_out[2][169]+ mul_add_t[2][169] + {4'b0000, e2[169]}%3329;
                                                                                                                                                                                     result[2][170] = decom_out[2][170]+ mul_add_t[2][170] + {4'b0000, e2[170]}%3329;
                                                                                                                                                                                     result[2][171] = decom_out[2][171]+ mul_add_t[2][171] + {4'b0000, e2[171]}%3329;
                                                                                                                                                                                     result[2][172] = decom_out[2][172]+ mul_add_t[2][172] + {4'b0000, e2[172]}%3329;
                                                                                                                                                                                     result[2][173] = decom_out[2][173]+ mul_add_t[2][173] + {4'b0000, e2[173]}%3329;
                                                                                                                                                                                     result[2][174] = decom_out[2][174]+ mul_add_t[2][174] + {4'b0000, e2[174]}%3329;
                                                                                                                                                                                     result[2][175] = decom_out[2][175]+ mul_add_t[2][175] + {4'b0000, e2[175]}%3329;
                                                                                                                                                                                     result[2][176] = decom_out[2][176]+ mul_add_t[2][176] + {4'b0000, e2[176]}%3329;
                                                                                                                                                                                     result[2][177] = decom_out[2][177]+ mul_add_t[2][177] + {4'b0000, e2[177]}%3329;
                                                                                                                                                                                     result[2][178] = decom_out[2][178]+ mul_add_t[2][178] + {4'b0000, e2[178]}%3329;
                                                                                                                                                                                     result[2][179] = decom_out[2][179]+ mul_add_t[2][179] + {4'b0000, e2[179]}%3329;
                                                                                                                                                                                     result[2][180] = decom_out[2][180]+ mul_add_t[2][180] + {4'b0000, e2[180]}%3329;
                                                                                                                                                                                     result[2][181] = decom_out[2][181]+ mul_add_t[2][181] + {4'b0000, e2[181]}%3329;
                                                                                                                                                                                     result[2][182] = decom_out[2][182]+ mul_add_t[2][182] + {4'b0000, e2[182]}%3329;
                                                                                                                                                                                     result[2][183] = decom_out[2][183]+ mul_add_t[2][183] + {4'b0000, e2[183]}%3329;
                                                                                                                                                                                     result[2][184] = decom_out[2][184]+ mul_add_t[2][184] + {4'b0000, e2[184]}%3329;
                                                                                                                                                                                     result[2][185] = decom_out[2][185]+ mul_add_t[2][185] + {4'b0000, e2[185]}%3329;
                                                                                                                                                                                     result[2][186] = decom_out[2][186]+ mul_add_t[2][186] + {4'b0000, e2[186]}%3329;
                                                                                                                                                                                     result[2][187] = decom_out[2][187]+ mul_add_t[2][187] + {4'b0000, e2[187]}%3329;
                                                                                                                                                                                     result[2][188] = decom_out[2][188]+ mul_add_t[2][188] + {4'b0000, e2[188]}%3329;
                                                                                                                                                                                     result[2][189] = decom_out[2][189]+ mul_add_t[2][189] + {4'b0000, e2[189]}%3329;
                                                                                                                                                                                     result[2][190] = decom_out[2][190]+ mul_add_t[2][190] + {4'b0000, e2[190]}%3329;
                                                                                                                                                                                     result[2][191] = decom_out[2][191]+ mul_add_t[2][191] + {4'b0000, e2[191]}%3329;
                                                                                                                                                                                     result[2][192] = decom_out[2][192]+ mul_add_t[2][192] + {4'b0000, e2[192]}%3329;
                                                                                                                                                                                     result[2][193] = decom_out[2][193]+ mul_add_t[2][193] + {4'b0000, e2[193]}%3329;
                                                                                                                                                                                     result[2][194] = decom_out[2][194]+ mul_add_t[2][194] + {4'b0000, e2[194]}%3329;
                                                                                                                                                                                     result[2][195] = decom_out[2][195]+ mul_add_t[2][195] + {4'b0000, e2[195]}%3329;
                                                                                                                                                                                     result[2][196] = decom_out[2][196]+ mul_add_t[2][196] + {4'b0000, e2[196]}%3329;
                                                                                                                                                                                     result[2][197] = decom_out[2][197]+ mul_add_t[2][197] + {4'b0000, e2[197]}%3329;
                                                                                                                                                                                     result[2][198] = decom_out[2][198]+ mul_add_t[2][198] + {4'b0000, e2[198]}%3329;
                                                                                                                                                                                     result[2][199] = decom_out[2][199]+ mul_add_t[2][199] + {4'b0000, e2[199]}%3329;
                                                                                                                                                                                     result[2][200] = decom_out[2][200]+ mul_add_t[2][200] + {4'b0000, e2[200]}%3329;
                                                                                                                                                                                     result[2][201] = decom_out[2][201]+ mul_add_t[2][201] + {4'b0000, e2[201]}%3329;
                                                                                                                                                                                     result[2][202] = decom_out[2][202]+ mul_add_t[2][202] + {4'b0000, e2[202]}%3329;
                                                                                                                                                                                     result[2][203] = decom_out[2][203]+ mul_add_t[2][203] + {4'b0000, e2[203]}%3329;
                                                                                                                                                                                     result[2][204] = decom_out[2][204]+ mul_add_t[2][204] + {4'b0000, e2[204]}%3329;
                                                                                                                                                                                     result[2][205] = decom_out[2][205]+ mul_add_t[2][205] + {4'b0000, e2[205]}%3329;
                                                                                                                                                                                     result[2][206] = decom_out[2][206]+ mul_add_t[2][206] + {4'b0000, e2[206]}%3329;
                                                                                                                                                                                     result[2][207] = decom_out[2][207]+ mul_add_t[2][207] + {4'b0000, e2[207]}%3329;
                                                                                                                                                                                     result[2][208] = decom_out[2][208]+ mul_add_t[2][208] + {4'b0000, e2[208]}%3329;
                                                                                                                                                                                     result[2][209] = decom_out[2][209]+ mul_add_t[2][209] + {4'b0000, e2[209]}%3329;
                                                                                                                                                                                     result[2][210] = decom_out[2][210]+ mul_add_t[2][210] + {4'b0000, e2[210]}%3329;
                                                                                                                                                                                     result[2][211] = decom_out[2][211]+ mul_add_t[2][211] + {4'b0000, e2[211]}%3329;
                                                                                                                                                                                     result[2][212] = decom_out[2][212]+ mul_add_t[2][212] + {4'b0000, e2[212]}%3329;
                                                                                                                                                                                     result[2][213] = decom_out[2][213]+ mul_add_t[2][213] + {4'b0000, e2[213]}%3329;
                                                                                                                                                                                     result[2][214] = decom_out[2][214]+ mul_add_t[2][214] + {4'b0000, e2[214]}%3329;
                                                                                                                                                                                     result[2][215] = decom_out[2][215]+ mul_add_t[2][215] + {4'b0000, e2[215]}%3329;
                                                                                                                                                                                     result[2][216] = decom_out[2][216]+ mul_add_t[2][216] + {4'b0000, e2[216]}%3329;
                                                                                                                                                                                     result[2][217] = decom_out[2][217]+ mul_add_t[2][217] + {4'b0000, e2[217]}%3329;
                                                                                                                                                                                     result[2][218] = decom_out[2][218]+ mul_add_t[2][218] + {4'b0000, e2[218]}%3329;
                                                                                                                                                                                     result[2][219] = decom_out[2][219]+ mul_add_t[2][219] + {4'b0000, e2[219]}%3329;
                                                                                                                                                                                     result[2][220] = decom_out[2][220]+ mul_add_t[2][220] + {4'b0000, e2[220]}%3329;
                                                                                                                                                                                     result[2][221] = decom_out[2][221]+ mul_add_t[2][221] + {4'b0000, e2[221]}%3329;
                                                                                                                                                                                     result[2][222] = decom_out[2][222]+ mul_add_t[2][222] + {4'b0000, e2[222]}%3329;
                                                                                                                                                                                     result[2][223] = decom_out[2][223]+ mul_add_t[2][223] + {4'b0000, e2[223]}%3329;
                                                                                                                                                                                     result[2][224] = decom_out[2][224]+ mul_add_t[2][224] + {4'b0000, e2[224]}%3329;
                                                                                                                                                                                     result[2][225] = decom_out[2][225]+ mul_add_t[2][225] + {4'b0000, e2[225]}%3329;
                                                                                                                                                                                     result[2][226] = decom_out[2][226]+ mul_add_t[2][226] + {4'b0000, e2[226]}%3329;
                                                                                                                                                                                     result[2][227] = decom_out[2][227]+ mul_add_t[2][227] + {4'b0000, e2[227]}%3329;
                                                                                                                                                                                     result[2][228] = decom_out[2][228]+ mul_add_t[2][228] + {4'b0000, e2[228]}%3329;
                                                                                                                                                                                     result[2][229] = decom_out[2][229]+ mul_add_t[2][229] + {4'b0000, e2[229]}%3329;
                                                                                                                                                                                     result[2][230] = decom_out[2][230]+ mul_add_t[2][230] + {4'b0000, e2[230]}%3329;
                                                                                                                                                                                     result[2][231] = decom_out[2][231]+ mul_add_t[2][231] + {4'b0000, e2[231]}%3329;
                                                                                                                                                                                     result[2][232] = decom_out[2][232]+ mul_add_t[2][232] + {4'b0000, e2[232]}%3329;
                                                                                                                                                                                     result[2][233] = decom_out[2][233]+ mul_add_t[2][233] + {4'b0000, e2[233]}%3329;
                                                                                                                                                                                     result[2][234] = decom_out[2][234]+ mul_add_t[2][234] + {4'b0000, e2[234]}%3329;
                                                                                                                                                                                     result[2][235] = decom_out[2][235]+ mul_add_t[2][235] + {4'b0000, e2[235]}%3329;
                                                                                                                                                                                     result[2][236] = decom_out[2][236]+ mul_add_t[2][236] + {4'b0000, e2[236]}%3329;
                                                                                                                                                                                     result[2][237] = decom_out[2][237]+ mul_add_t[2][237] + {4'b0000, e2[237]}%3329;
                                                                                                                                                                                     result[2][238] = decom_out[2][238]+ mul_add_t[2][238] + {4'b0000, e2[238]}%3329;
                                                                                                                                                                                     result[2][239] = decom_out[2][239]+ mul_add_t[2][239] + {4'b0000, e2[239]}%3329;
                                                                                                                                                                                     result[2][240] = decom_out[2][240]+ mul_add_t[2][240] + {4'b0000, e2[240]}%3329;
                                                                                                                                                                                     result[2][241] = decom_out[2][241]+ mul_add_t[2][241] + {4'b0000, e2[241]}%3329;
                                                                                                                                                                                     result[2][242] = decom_out[2][242]+ mul_add_t[2][242] + {4'b0000, e2[242]}%3329;
                                                                                                                                                                                     result[2][243] = decom_out[2][243]+ mul_add_t[2][243] + {4'b0000, e2[243]}%3329;
                                                                                                                                                                                     result[2][244] = decom_out[2][244]+ mul_add_t[2][244] + {4'b0000, e2[244]}%3329;
                                                                                                                                                                                     result[2][245] = decom_out[2][245]+ mul_add_t[2][245] + {4'b0000, e2[245]}%3329;
                                                                                                                                                                                     result[2][246] = decom_out[2][246]+ mul_add_t[2][246] + {4'b0000, e2[246]}%3329;
                                                                                                                                                                                     result[2][247] = decom_out[2][247]+ mul_add_t[2][247] + {4'b0000, e2[247]}%3329;
                                                                                                                                                                                     result[2][248] = decom_out[2][248]+ mul_add_t[2][248] + {4'b0000, e2[248]}%3329;
                                                                                                                                                                                     result[2][249] = decom_out[2][249]+ mul_add_t[2][249] + {4'b0000, e2[249]}%3329;
                                                                                                                                                                                     result[2][250] = decom_out[2][250]+ mul_add_t[2][250] + {4'b0000, e2[250]}%3329;
                                                                                                                                                                                     result[2][251] = decom_out[2][251]+ mul_add_t[2][251] + {4'b0000, e2[251]}%3329;
                                                                                                                                                                                     result[2][252] = decom_out[2][252]+ mul_add_t[2][252] + {4'b0000, e2[252]}%3329;
                                                                                                                                                                                     result[2][253] = decom_out[2][253]+ mul_add_t[2][253] + {4'b0000, e2[253]}%3329;
                                                                                                                                                                                     result[2][254] = decom_out[2][254]+ mul_add_t[2][254] + {4'b0000, e2[254]}%3329;
                                                                                                                                                                                     result[2][255] = decom_out[2][255]+ mul_add_t[2][255] + {4'b0000, e2[255]}%3329;
                                                                                                                                                                                    
                                           
                                                                                                                                                  end
                                                                                                                                                  end
                                                                                                                                              
                                                                                                                                              
                                           
                                                                    
                                                      end
                                                      end       
                                       
                                    
                                   
                          endmodule