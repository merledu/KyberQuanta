`timescale 1ns / 1ps

module tb_encode;

    // Parameters
    parameter D = 12;
    parameter BYTE_LEN = 32;
    parameter NUM_INPUTS = 256;

    // DUT inputs and outputs
    logic signed [15:0] F [NUM_INPUTS-1:0]; // Input 16-bit signed array
    logic [7:0] B [BYTE_LEN * D - 1:0];    // Output byte array

    // Instantiate the DUT
    encode #(
        .D(D),
        .BYTE_LEN(BYTE_LEN)
    ) dut (
        .F(F),
        .B(B)
    );

    // Testbench variables
    integer i;

    initial begin
        // Initialize the input array F
        F= '{106, 1613, 2786, 3016, 2498, 120, 3302, 224, 2957, 1447, 625, 2861, 1413, 594, 2556, 129, 1845, 1880, 1991, 2996, 1764, 2200, 381, 714, 1712, 2111, 457, 481, 1395, 3282, 2773, 1311, 2592, 3083, 2877, 644, 1347, 401, 1985, 1947, 3079, 1863, 623, 1743, 1337, 3239, 763, 2844, 2047, 1084, 2264, 1763, 3082, 676, 2004, 2235, 2468, 2135, 2921, 1036, 2271, 2854, 1549, 1986, 717, 913, 2686, 2405, 1016, 498, 2740, 1523, 1066, 1448, 3004, 2242, 2793, 2467, 2459, 2121, 2917, 648, 2053, 1142, 1564, 1344, 777, 2276, 153, 760, 1048, 1487, 1425, 2278, 430, 1655, 2265, 2123, 3202, 756, 611, 970, 2760, 1761, 1039, 1288, 1487, 1874, 797, 1934, 3060, 468, 3122, 1833, 1114, 3007, 1971, 1476, 12, 1569, 487, 1258, 3279, 3092, 2406, 2470, 2751, 866, 2719, 873, 1353, 2423, 443, 1985, 1403, 1164, 599, 580, 1098, 2400, 726, 2503, 2431, 288, 1939, 1330, 1806, 562, 632, 2591, 2450, 1209, 2977, 2657, 884, 548, 2837, 2847, 988, 2846, 1935, 552, 2576, 1309, 1308, 1122, 1947, 2606, 1889, 345, 144, 869, 147, 2170, 468, 2580, 609, 2887, 1610, 464, 2806, 222, 45, 2483, 3318, 584, 758, 1348, 2968, 606, 210, 286, 653, 1826, 1437, 1264, 1016, 1182, 1847, 2778, 2134, 1656, 644, 1982, 0, 453, 174, 1489, 1960, 1905, 1567, 621, 2490, 1780, 1490, 3123, 2322, 1239, 923, 51, 2573, 1854, 1480, 848, 1909, 2361, 1365, 380, 1553, 2868, 88, 2184, 428, 1367, 766, 3103, 2570, 473, 223, 2391, 464, 1624, 1161, 755, 229, 437, 2876, 2306, 1658, 1490, 2722, 2955, 676, 2005, 1197, 1817};

        // Wait for the combinational logic to propagate
        #10;

        // Display the encoded output byte array
        $display("Encoded byte array B:");
        for (i = 0; i < BYTE_LEN * D; i = i + 1) begin
            $display("B[%0d] = %0d", i, B[i]);
        end

        // Finish simulation
        $finish;
    end

endmodule
