`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/24/2025 10:55:23 PM
// Design Name: 
// Module Name: KPKE_decrypt_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////




module KPKE_decrypt_tb;

    // Parameters (must match the DUT)
    localparam DK_BYTES  = 1152;
    localparam C_BYTES   = 1088;
    localparam MSG_BYTES = 32;

    // DUT signals
    logic clk;
    logic rst;
    logic start;
    logic [7:0] dk_PKE [0:DK_BYTES-1];
    logic [7:0] c      [0:C_BYTES-1];
    logic done_1;
    logic [7:0] m      [0:MSG_BYTES-1];
    logic done_encode_debug;

    // Instantiate the DUT
    K_PKE_Decrypt #(
        .DK_BYTES(DK_BYTES),
        .C_BYTES(C_BYTES),
        .MSG_BYTES(MSG_BYTES)
    ) dut (
        .clk(clk),
        .rst(rst),
        .start(start),
        .dk_PKE(dk_PKE),
        .c(c),
        .done_1(done_1),
        .m(m),
        .done_encode_debug(done_encode_debug)
    );

    // Clock generation: 100 MHz
    initial clk = 0;
    always #5 clk = ~clk;

    // Test stimulus
    reg [9215:0] dk_PKE_bits;
    reg [8703:0] c_bits;

    initial begin
        integer i;

        // Initial conditions
        rst   = 1;
        start = 0;

        // Assign packed test vectors
     dk_PKE_bits = 9216'h125C69B3959521000369BA3470AB58AC1CEE7D108A48F619CB90D35F507E07201A72B315BB3C613F55BF9EE231C2D29ACFD0727F530A7CCBD96EF8BB56A01BB5970C8127FF465565C76C509C629E29E5D080056CB3D854132AC2BAC46A9F56203257A825BC10C8CCD083917672961FAD2B47405C67B06B7733E6F08201D513AABD5A002057F5BD3C47BA51177892C7E831A01691342E43648A138B03A80BADC6DA993E761C4A69037B2AAA4910FC844247CBE50F71741525D056480B96ABF003C5570A5CB99A0E57432E8B1B491A00A1CA63891B94CFD7345E941D680626BA241730650678347B5540A8B9322B1321A8C8F7E1849A2EB0DC4442CAF938405DCA74A3A820F333A60070D65368209429780B29F691B7E4D34F15944EEACB422C1247464B3A945424BCA214B11E28E415B078F13B067EB62496B5F858B0E42CA006410388CA5245EF1D25BE1AD99054A5D4BA701992F4BE2710A49A92E28936B62799A12A584991AADF5724CA462913415B0998BB571838059624C9BDE4AD6314AA34230ACF59A495E5D11AAB992FC7D40E2371B3338426D79557B8C10AB5670788768BA5CB81B32C8865D534912554644164B55F9F6316ADD5F11579AC9E90D64F33F14D503BCC62200777AD690695313CAB453A3E72796AB4E3BF983BDA3AA0F03E059527D3A662D66C4B006AA3EC69CCB0C79AE0AEB4C995AFD34F0685BBB495A6893C0BCE41FDA81B1949375A11995DAFD4BC6159C73006B01A81AF4D46F443A246963AE4499B9245B0DA7413221901F934038FC279793811418F13C93879C12FF9C3817A592923022C466053F631030AE01CC5F3AB1265C8851ABDD6CB3D3A3FA7E66E5835D700200239020B0F51F380D92C0F7B59211A79CDD0C90CF29252F5B3451071A02496AEFA7F45D2F29355954B3AF0A156299EF5D3B498E66CB5E39C106391B29C598C074A2927302A330435644D43E564992F77337DC6C36147977A016B137B44B06DD5EB5C98C6AE573C66A94C13633A2DBCE151F88B8BDA291B452717AB9EB6A7BF3124DF8926A9315B4280E33961B8890166AD513B7CA57AEE03F9CC92023CA85765460B8AAF85F476EB057689CF0CB877BDE4345706C82AF66CB14853AE75928B27D265AAD0B945E77583B71A47CD523CEF6CE6F92EFA3435878B3FB48A55EAEB8A326CA8912C214AC794A2C54F778C9F630C098B38AFF8725C007F9823421597944611B8840B921A6A10CB23F41FE9099B99C613D22C6AB9419A58F211902F4251E56A852B3AC0940FFA6E70053DB6E634B5E6F63366A15239A0B347CF8C33EDB9B35F0B12BE62E9EB5786101AA819B547EF2B765F2E381A2884F262471B90023856C4CD266B351B30A4A2B2FABFB234AB7A836C968C1B32860C521535875F295AD9A0FB992BF90C1B5B18CC27910C1C40A501B053B270B20586B4F70864217DBE6C7F4E4BF4A938FF0531497D05F5B6E668BA84BA495A8A84D89EA2C1FA0CEB1412753FCBFCBC9B9BC7A0AA3A22D5B310437A185058A0B0451892F6C3A644028600029CA1B33C535922F4BCA46B20321CA305224787CB73178E2AD2C0A9921C93E81DB8027559747542F5707E2B71AC72E607F79B855634;
     c_bits = 8704'hC6D205D9AF4FE4A3120F3331751C279915D9C34CC3FE10C0C8B60B258D1ACB60C6D47B238FF4390E9AACC3C5CE4CF5BBC6CEA9550B65656753C1EC9E13DC3F5FF0A641B8727D4CE1918530F76806CC839D0D337E6E621E222B0CE43B6E2B0E1FD94882B4ACB9FBB1202271700FDE7CDF79C8B62893F71C270F63DF36C384FD10C188EC71BABAE659D1180A793C9FAC6AC9E07BB32AB07FBED6517FBE5EAD3027438387E60E38DACB769523417A7A7C21EB94B028AEC115EA145664E56C57C454774F1B7E45A20A2B6C7599B1D89878802837C7F7B116A0F6B29668CA764033E9CB17F17C24F5CD6B69FE6814DA94AFCB24FB1614C35CCA90EAE20BE29C7886FEEDC60E7DAB55360890F372869A1DE7916C9004642B47BEE53BEA161477F2F560ED88E0C6C36F39E8FC60655E499DB16B7DDA4B23A6017CD7E750E5A345B7DA4233938DFD39D4A189275A60C322ED6A0187EAAF9A857CFA76AC820107BC6F280C7B6025BA092BE89204F9860DB796E3114B68396B1FDF001629FFDB3FEB7E90AA70329D9FA91430A1DD6248F601A52A2E0A9397172365D40E200300BC0A047420A6185D1C0649DAE724000C720F70D0D6E982E8C8AF8BE70194FE06B889142444E7B9E8F347496A04EFD3BAECD09549A55FE1F4B4888E4B817E7C0E780D9FF0EA888ED99CF99A157E9A11964AB75D2AB395EEAB034B8C60BEC94A5D61258598EFA2146820D908E76EA1FD6B626DCEA8EC7F4CFAFF7DF3FB2EFBF8C1CEDB4DEC9B4A1FF31FF61987D20B155220CD1934A4010CB703C98D3BD66123E6DD6CE178BCF43AA189952F5FB193E383FF4A270FEF8C7CE1F7606090FBFB7195CC5708F841CC8CD0C5F4DB4C31D74674198F4A20E2EF57CD3573BB3C68CEB081F7E38E65A898524BDEBE8A3E5E729D8BACFC29C79E8160D55C9BDD299E30BA85FB5CD49FD3033CBB2E741F0B9138824699BC4316CF4B93A2119DBD68954570A0CD9CD6561963CFDA8AE7C7B5EF07AB3D158AF58D638019E0D1AC9514CD5782F30A782259E2E314270F463A801EA2E7293136633F2D9AB2D7E973961514367D6B701CFDD4CC2C29762AACBD1A9755C9683885C4EF4FC5E775F7FE0D1C674AB552D554FFCA1B68B052818C27CB14A2224EC145B16CE02DE211015D3A1A09603A519C0678E4FD2ACF7900C977A99B751458EBCD98D6B85DEEE5E99BE9DCA09BEDA2C41C59079E05B32207095117D1F78CA784391D5717B340DFA9C00D473896C0EF572A94047D64A5D3ECF874F826A8B34E31D516A6F374FEE337FF843980AC884FB0FAB2B498F593AB51B977A8AF4AB0F866EFA893B3C649077B30EB0D682E24FB2126268C3F910FED392DF5E079D2121AA70CEE9135C2C8346CF370EF42093719BC219564709B614946A12A63B2943AD483E1F74B04AE2E071904C9C7BB5B0E11F87B08009DE27E359DEB77EB14F462CED4887D75C3555A231EA282B217D74AFE4177D80F73C1BAEAA66F288D1CE9FC91F9FE6B87CF6ED5E0F750DE9DB820B4632AD7B9A6DF;
            
             
        // Bit-slice into byte arrays
        for (i = 0; i < DK_BYTES; i = i + 1)
            dk_PKE[i] = dk_PKE_bits[8*(DK_BYTES - i) - 1 -: 8];

        for (i = 0; i < C_BYTES; i = i + 1)
            c[i] = c_bits[8*(C_BYTES - i) - 1 -: 8];

        // Reset sequence
        #5000;
        rst = 0;
        

        // Start signal pulse
        start = 1;
        #400000;
        

        // Wait for decryption to finish
        wait (done_1);

        // Display decrypted message
        $display("Decryption complete. Output message:");
        for (i = 0; i < MSG_BYTES; i = i + 1)
            $write("%02x ", m[i]);
        $display();

        #20;
        $finish;
    end

endmodule
