`timescale 1ns / 1ps
module encryption #( 
    parameter k = 3,
    parameter ELL = 16,
    parameter NUM_COEFFS = 256,
    parameter Q = 3329
)(
  input logic clk,
  input logic rst,
  input logic [7:0] pk[1183:0],    
  input logic [7:0] mess [32-1:0], 
  input [255:0] r,     
  output logic [15:0] A [0:2][0:2][0:255],
  output logic [ 16-1:0] T_hat_0 [0:256-1],
  output logic [ 16-1:0] T_hat_1 [0:256-1],
  output logic [ 16-1:0] T_hat_2 [0:256-1],
  output logic [ 16-1:0] m_dec [0:256-1],
  output logic [255:0] rho_t,
  output logic [11:0] y [0:2][255:0],
  output logic [11:0] e1 [0:2][255:0],
  output logic [15:0] y_ntt [0:2][255:0],
  output logic start_ntt,
  output logic start_inverse,
  output logic [15:0] mult_out_00 [255:0],
  output logic [15:0] mult_out_01 [255:0],
  output logic [15:0] mult_out_02 [255:0],
  output logic [15:0] mult_out_10 [255:0],
  output logic [15:0] mult_out_11 [255:0],
  output logic [15:0] mult_out_12 [255:0],
  output logic [15:0] mult_out_20 [255:0],
  output logic [15:0] mult_out_21 [255:0],
      output logic [15:0] mult_out_22 [255:0],
      output logic  done9_mul,
      output logic  done10_mul,
      output logic  done11_mul,
      output logic [15:0] mult_out_1 [255:0],
      output logic [15:0] mult_out_2 [255:0],
      output logic [15:0] mult_out_3 [255:0],
       output logic done0_mul,
        output logic  done1_mul,
       output  logic  done2_mul,
       output  logic  done3_mul,
       output  logic  done4_mul,
       output  logic  done5_mul,
       output  logic  done6_mul,
        output logic done7_mul,
        output logic  done8_mul,
        output logic start_mul, 
        output logic [15:0] mul_add [0:2][255:0],          
         output   logic  done0_ntt,
          output  logic done1_ntt,
         output   logic done2_ntt,
            output logic done10_ntt,
               output logic done11_ntt,
               output logic done12_ntt,
               output logic [31:0] in_1 [256-1:0],
                 output logic [31:0] in_2 [256-1:0],
                 output logic [31:0] in_3 [256-1:0],
                 output logic [31:0] in_4 [256-1:0],
               output logic [31:0] in_5 [256-1:0],
           output logic [31:0] in_6 [256-1:0], 
           output logic  [15:0] decom_out [0:256-1],
           output logic [11:0] e2 [255:0],
           output logic [31:0] v [255:0],
            output logic done13_ntt,
           output logic done14_ntt,
            output logic done15_ntt,
                 output logic [31:0] u [0:2][255:0] , 
                 output logic [15:0] mul_add_t[0:2][255:0], 
                 output logic [15:0] com_out [0:2][255:0],
                 output logic [15:0] comp_v [255:0], 
                 output logic [7:0] encode_u [0:2] [256-1:0],
                 output logic [7:0] encode_v  [255:0]

      );
    

    logic [7:0] pk_slice0 [0:383];
    logic [7:0] pk_slice1 [0:383];
    logic [7:0] pk_slice2 [0:383];
    logic  done9_shake, done10_shake, done11_shake, done12_shake, done13_shake, done14_shake,done15_shake;
    logic  done0_cbd, done1_cbd, done2_cbd, done3_cbd, done4_cbd, done5_cbd,done6_cbd;
    logic [7:0] parse_array1 [767:0];
    logic [7:0] parse_array2 [767:0];
    logic [7:0] parse_array3 [767:0];
    logic [7:0] parse_array4 [767:0];
    logic [7:0] parse_array5 [767:0];
    logic [7:0] parse_array6 [767:0];
    logic [7:0] parse_array7 [767:0];
    logic [7:0] parse_array8 [767:0];
    logic [7:0] parse_array9 [767:0];
    logic start1;
    logic done0, done1, done2, done3, done4, done5, done6, done7, done8, done9;
    logic done0_shake,done1_shake,done2_shake,done3_shake,done4_shake,done5_shake,done6_shake,done7_shake,done8_shake;
    logic all_shake_done;
    logic [7:0] prf_bytes_0 [127:0];
    logic [7:0] prf_bytes_1 [127:0];
    logic [7:0] prf_bytes_2 [127:0];
    logic [7:0] prf_bytes_3 [127:0];
    logic [7:0] prf_bytes_4 [127:0];
    logic [7:0] prf_bytes_5 [127:0];
    logic [7:0] prf_bytes_6 [127:0];
    logic [1023:0] prf_0, prf_1, prf_2, prf_3, prf_4, prf_5, prf_6;
    logic  start_parse, start_cbd, start_prf;
    logic [15:0] zetas [127:0];
    logic ntt_started;
    logic mul;
    logic [268-1:0] r0;
    logic [268-1:0] r1;
    logic [268-1:0] r2;
    logic [268-1:0] r3;
    logic [268-1:0] r4;
    logic [268-1:0] r5;
   

    
    
    assign pk_slice0 = pk[383:0];
    assign pk_slice1 = pk[767:384];
    assign pk_slice2 = pk[1151:768];
   
assign rho_t = {
           pk[1152], pk[1153], pk[1154], pk[1155],
           pk[1156], pk[1157], pk[1158], pk[1159],
           pk[1160], pk[1161], pk[1162], pk[1163],
           pk[1164], pk[1165], pk[1166], pk[1167],
           pk[1168], pk[1169], pk[1170], pk[1171],
           pk[1172], pk[1173], pk[1174], pk[1175],
           pk[1176], pk[1177], pk[1178], pk[1179],
           pk[1180], pk[1181], pk[1182], pk[1183]
       };


    decode #(.ELL(16), .NUM_COEFFS(256), .BYTE_COUNT(384)) dec0 (
        .byte_array(pk_slice0),
        .len(384),
        .coeffs(T_hat_0)
    );

    decode #(.ELL(16), .NUM_COEFFS(256), .BYTE_COUNT(384)) dec1 (
        .byte_array(pk_slice1),
        .len(384),
        .coeffs(T_hat_1)
    );

    decode #(.ELL(16), .NUM_COEFFS(256), .BYTE_COUNT(384)) dec2 (
        .byte_array(pk_slice2),
        .len(384),
        .coeffs(T_hat_2)
    );
   logic [7:0] mess [32-1:0];
    assign mess[0]  = 8'hEB;
   assign mess[1]  = 8'h4A;
   assign mess[2]  = 8'h7C;
   assign mess[3]  = 8'h66;
   assign mess[4]  = 8'hEF;
   assign mess[5]  = 8'h4E;
   assign mess[6]  = 8'hBA;
   assign mess[7]  = 8'h2D;
   assign mess[8]  = 8'hDB;
   assign mess[9]  = 8'h38;
   assign mess[10] = 8'hC8;
   assign mess[11] = 8'h8D;
   assign mess[12] = 8'h8B;
   assign mess[13] = 8'hC7;
   assign mess[14] = 8'h06;
   assign mess[15] = 8'hB1;
   assign mess[16] = 8'hD6;
   assign mess[17] = 8'h39;
   assign mess[18] = 8'h00;
   assign mess[19] = 8'h21;
   assign mess[20] = 8'h98;
   assign mess[21] = 8'h17;
   assign mess[22] = 8'h2A;
   assign mess[23] = 8'h7B;
   assign mess[24] = 8'h19;
   assign mess[25] = 8'h42;
   assign mess[26] = 8'hEC;
   assign mess[27] = 8'hA8;
   assign mess[28] = 8'hF6;
   assign mess[29] = 8'hC0;
   assign mess[30] = 8'h01;
   assign mess[31] = 8'hBA;

  decode #(.ELL(16), .NUM_COEFFS(256),.BYTE_COUNT(32)) dec4 (
                         .byte_array(mess),
                         .len(32),
                         .coeffs(m_dec)
                     );     
              //--------------------------XOF 1--------------------------------------
    logic [276-1:0] datain;
    logic [6144-1:0] xof;
    
   assign datain = {4'hF,8'h00, 8'h00,rho_t};
   assign message = datain; 
//   assign done0_shake = 1'b1;
    sponge #(
     .msg_len(276),
     .d_len(6144),
     .capacity(256),
     .r(1600 - 256)
 ) shake1(
        .clk(clk),
        .reset(rst),
        .start(start1),
        .message(datain),
        .z(xof),
        .done(done0_shake)
    );
            
           
           //--------------------------XOF 2--------------------------------------
              logic [276-1:0] datain2;
                   logic [6144-1:0] xof2;
//                  assign message = datain2; 
                   assign datain2 = {4'hF ,8'h00, 8'h02,rho_t};     
                    
                   sponge #(
                    .msg_len(276),
                    .d_len(6144),
                    .capacity(256),
                    .r(1600 - 256)
                ) shake2(
                       .clk(clk),
                       .reset(rst),
                       .start(start1),
                       .message(datain2),
                       .z(xof2),
                       .done(done1_shake)
                   ); 
                    
                 //--------------------------XOF 3--------------------------------------
               logic [276-1:0] datain3;
               logic [6144-1:0] xof3;
//                        assign message = datain3;                           
               assign datain3 = {4'hF , 8'h00, 8'h11,rho_t };      
               sponge #(
                    .msg_len(276),
                     .d_len(6144),
                     .capacity(256),
                     .r(1600 - 256)
                                  ) shake3(
                                        .clk(clk),
                                         .reset(rst),
                                         .start(start1),
                                        .message(datain3),
                                          .z(xof3),
                                           .done(done2_shake)
                                                  );
   
                    // --------------------------XOF 4--------------------------------------
              logic [276-1:0] datain4;
              logic [6144-1:0] xof4;
//                                                            assign message = datain4; 
              assign datain4 = {4'hF ,  8'h01 , 8'h00,rho_t };
              sponge #(
                        .msg_len(276),
                         .d_len(6144),
                         .capacity(256),
                         .r(1600 - 256)
                   ) shake4 (
                              .clk(clk),
                             .reset(rst),
                             .start(start1),
                            .message(datain4),
                             .z(xof4),
                             .done( done3_shake)
                                        );        
                  
                    // --------------------------XOF 5--------------------------------------
                         logic [276-1:0] datain5;
                  logic [6144-1:0] xof5;
//                assign message = datain5; 
            assign datain5 = {4'hF ,  8'h01 , 8'h01,rho_t };
        sponge #(
                      .msg_len(276),
                      .d_len(6144),
                      .capacity(256),
                       .r(1600 - 256)
                                       )
                 shake5 (
                         .clk(clk),
                         .reset(rst),
                         .start(start1),
                         .message(datain5),
                         .z(xof5),
                         .done( done4_shake)
                          );  
                 
                    // --------------------------XOF 6--------------------------------------
                       logic [276-1:0] datain6;
                       logic [6144-1:0] xof6;
//                       assign message = datain6; 
                       assign datain6 = {4'hF ,  8'h1 , 8'h2,rho_t };
                       sponge #(
                       .msg_len(276),
                       .d_len(6144),
                       .capacity(256),
                       .r(1600 - 256)
                       ) shake6 (
                       .clk(clk),
                        .reset(rst),
                        .start(start1),
                        .message(datain6),
                        .z(xof6),
                        .done( done5_shake)
                        );
                  
               // --------------------------XOF 7--------------------------------------
                   logic [276-1:0] datain7;
                   logic [6144-1:0] xof7;
//                    assign message = datain7; 
                   assign datain7 = {4'hF ,  8'h02 , 8'h00,rho_t };
                   sponge #(
                   .msg_len(276),
                   .d_len(6144),
                   .capacity(256),
                   .r(1600 - 256)
                   ) shake7 (
                   .clk(clk),
                   .reset(rst),
                   .start(start1),
                   .message(datain7),
                   .z(xof7),
                   .done( done6_shake)
                    );
   
                    // --------------------------XOF 8--------------------------------------
                     logic [276-1:0] datain8;
                     logic [6144-1:0] xof8;
//                     assign message = datain8; 
                     assign datain8 = {4'hF ,  8'h02 , 8'h01,rho_t };
                      sponge #(
                       .msg_len(276),
                       .d_len(6144),
                       .capacity(256),
                        .r(1600 - 256)
                         ) shake8 (
                          .clk(clk),
                           .reset(rst),
                            .start(start1),
                            .message(datain8),
                            .z(xof8),
                             .done( done7_shake)
                              );
                                                                                                          
                                                                                                          // --------------------------XOF 9--------------------------------------
          logic [276-1:0] datain9;
          logic [6144-1:0] xof9;
//        assign message = datain9; 
          assign datain9 = {4'hF ,  8'h2 , 8'h2,rho_t };
          sponge #(
           .msg_len(276),
           .d_len(6144),
           .capacity(256),
           .r(1600 - 256)
            ) shake9 (
            .clk(clk),
            .reset(rst),
            .start(start1),
            .message(datain9),
            .z(xof9),
            .done( done8_shake)
             );
       parse parse_00 (.clk(clk),.rst(rst),.start(done0_shake),.done(done0), .B(parse_array1), .a(A[0][0]));
       parse parse_01 (.clk(clk),.rst(rst),.start(done1_shake),.done(done1),.B(parse_array2), .a(A[0][1]));
       parse parse_02 (.clk(clk),.rst(rst),.start(done2_shake),.done(done2),.B(parse_array3), .a(A[0][2]));
       
       parse parse_10 (.clk(clk),.rst(rst),.start(done3_shake),.done(done3),.B(parse_array4), .a(A[1][0]));
       parse parse_11 (.clk(clk),.rst(rst),.start(done4_shake),.done(done4),.B(parse_array5), .a(A[1][1]));
       parse parse_12 (.clk(clk),.rst(rst),.start(done4_shake),.done(done5),.B(parse_array6), .a(A[1][2]));
       
       parse parse_20 (.clk(clk),.rst(rst),.start(done4_shake),.done(done6),.B(parse_array7), .a(A[2][0]));
       parse parse_21 (.clk(clk),.rst(rst),.start(done4_shake),.done(done7),.B(parse_array8), .a(A[2][1]));
       parse parse_22 (.clk(clk),.rst(rst),.start(done8_shake),.done(done8),.B(parse_array9), .a(A[2][2]));
       

     
//     //-----------------prf0-------------------------
    
     
     assign r0 = {4'h1111, 8'h00,r}; 
     assign r1 = {4'h1111, 8'h01,r};
      assign r2 = {4'h1111, 8'h02,r};
         assign r3 = {4'h1111, 8'h03,r};  
            assign r4 = {4'h1111, 8'h04,r}; 
             assign r5 = {4'h1111, 8'h05,r};
             
     sponge #(.msg_len(268),
      .d_len(1024), 
      .capacity(512),
       .r(1600 - 512))
        prf0 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r0),
         .z(prf_0),
         .done(done9_shake)
     );
     
  
     sponge #(.msg_len(268), 
     .d_len(1024), 
     .capacity(512), 
     .r(1600 - 512)) 
     prf1 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r1),
         .z(prf_1),
         .done(done10_shake)
     );
     
    
     sponge #(.msg_len(268), 
     .d_len(1024), 
     .capacity(512),
      .r(1600 - 512)) 
      prf2 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r2),
         .z(prf_2),
         .done(done11_shake)
     );
   
  
     sponge #(.msg_len(268),
      .d_len(1024), 
      .capacity(512),
       .r(1600 - 512))
        prf3 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r3),
         .z(prf_3),
         .done(done12_shake)
     );
     
   
     sponge #(.msg_len(268),
      .d_len(1024),
       .capacity(512),
        .r(1600 - 512)) 
        prf4 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r4),
         .z(prf_4),
         .done(done13_shake)
     );
     
     
    
     sponge #(.msg_len(268),
      .d_len(1024),
       .capacity(512),
        .r(1600 - 512))
      prf5 (
         .clk(clk),
         .reset(rst),
         .start(done8),
         .message(r5),
         .z(prf_5),
         .done(done14_shake)
     );
                  
        CBD cbd0 (.clk(clk), .reset(rst), .start(done14_shake), .done(done0_cbd), .byte_array(prf_bytes_0), .len(128), .f(y[0]));
        CBD cbd1 (.clk(clk), .reset(rst), .start(done14_shake), .done(done1_cbd), .byte_array(prf_bytes_1), .len(128), .f(y[1]));
        CBD cbd2 (.clk(clk), .reset(rst), .start(done14_shake), .done(done2_cbd), .byte_array(prf_bytes_2), .len(128), .f(y[2]));
        
        CBD cbd3 (.clk(clk), .reset(rst), .start(done14_shake), .done(done3_cbd), .byte_array(prf_bytes_3), .len(128), .f(e1[0]));
        CBD cbd4 (.clk(clk), .reset(rst), .start(done14_shake), .done(done4_cbd), .byte_array(prf_bytes_4), .len(128), .f(e1[1]));
        CBD cbd5 (.clk(clk), .reset(rst), .start(done14_shake), .done(done5_cbd), .byte_array(prf_bytes_5), .len(128), .f(e1[2]));
        

        logic [268-1:0] r6;
        assign r6 = {4'h1111, 8'h06,r}; 
        sponge #(.msg_len(268),
             .d_len(1024), 
             .capacity(512),
              .r(1600 - 512))
               prf6 (
                .clk(clk),
                .reset(rst),
                .start(done8),
                .message(r6),
                .z(prf_6),
                .done(done15_shake)
            );
               CBD cbd6  (
                  .clk(clk), 
                           .reset(rst), 
                           .start(done14_shake), 
                           .done(done6_cbd), 
                           .byte_array(prf_bytes_6), 
                           .len(128), 
                           .f(e2)
              );
              
               assign start_ntt = (done5_cbd && !done0_ntt && !done1_ntt && !done2_ntt);
               
                   ntt ntt_y0 (.clk(clk), .reset(rst), .f(y[0]), .start(start_ntt), .done(done0_ntt), .f_hat(y_ntt[0]));
                   ntt ntt_y1 (.clk(clk), .reset(rst), .f(y[1]), .start(start_ntt), .done(done1_ntt),.f_hat(y_ntt[1]));
                   ntt ntt_y2 (.clk(clk), .reset(rst), .f(y[2]), .start(start_ntt), .done(done2_ntt),.f_hat(y_ntt[2]));
           
                      
                     assign start_mul = (done0_ntt && done1_ntt && done2_ntt);
                  
                      multiply_ntts mul_00 (.clk(clk), .reset(rst),.f(A[0][0]), .g(y_ntt[0]), .zetas(zetas), .h(mult_out_00), .start(start_mul), .done(done0_mul));
                      multiply_ntts mul_01 (.clk(clk), .reset(rst),.f(A[0][1]), .g(y_ntt[1]), .zetas(zetas), .h(mult_out_01),.start(start_mul), .done(done1_mul));
                      multiply_ntts mul_02 (.clk(clk), .reset(rst),.f(A[0][2]), .g(y_ntt[2]), .zetas(zetas), .h(mult_out_02),.start(start_mul), .done(done2_mul));
                  
                      multiply_ntts mul_10 (.clk(clk), .reset(rst),.f(A[1][0]), .g(y_ntt[0]), .zetas(zetas), .h(mult_out_10), .start(start_mul), .done(done3_mul));
                      multiply_ntts mul_11 (.clk(clk), .reset(rst),.f(A[1][1]), .g(y_ntt[1]),.zetas(zetas), .h(mult_out_11), .start(start_mul), .done(done4_mul));
                      multiply_ntts mul_12 (.clk(clk), .reset(rst),.f(A[1][2]), .g(y_ntt[2]), .zetas(zetas),.h(mult_out_12), .start(start_mul), .done(done5_mul));
                  
                      multiply_ntts mul_20 (.clk(clk), .reset(rst),.f(A[2][0]), .g(y_ntt[0]),.zetas(zetas), .h(mult_out_20), .start(start_mul),.done(done6_mul));
                      multiply_ntts mul_21 (.clk(clk), .reset(rst),.f(A[2][1]), .g(y_ntt[1]), .zetas(zetas),.h(mult_out_21), .start(start_mul), .done(done7_mul));
                      multiply_ntts mul_22 (.clk(clk), .reset(rst),.f(A[2][2]), .g(y_ntt[2]), .zetas(zetas),.h(mult_out_22), .start(start_mul), .done(done8_mul));

                      
                      multiply_ntts
                          mult_1 (
                              .clk(clk),
                              .reset(rst),
                              .f(T_hat_0),  // T_hat_0_16 is a 16-bit array
                              .g(y_ntt[0]),  // y_ntt_0_16 is now a 1D array
                              .zetas(zetas),
                              .h(mult_out_1),
                              .start(start_mul),
                              .done(done9_mul)
                          );
                      
                      multiply_ntts
                          mult_2 (
                              .clk(clk),
                              .reset(rst),
                              .f(T_hat_1),  // T_hat_1_16 is a 16-bit array
                              .g(y_ntt[1]),  // y_ntt_1_16 is now a 1D array
                              .zetas(zetas),
                              .h(mult_out_2),
                              .start(start_mul),
                              .done(done10_mul)
                          );
                      
                      multiply_ntts
                          mult_3 (
                              .clk(clk),
                              .reset(rst),
                              .f(T_hat_2),  
                              .g(y_ntt[2]),  
                              .zetas(zetas),
                              .h(mult_out_3),
                              .start(start_mul),
                              .done(done11_mul)
                          );
                          assign start_inverse = (done3_mul && done4_mul && done5_mul );
                          
                          ////AT x Y inverse
//                          logic  [31:0] in_1 [256-1:0];
                          
                          inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_1 (
                              .clk(clk),
                              .rst(rst),
                              .f(mul_add[0]),
                              .start_ntt(start_inverse),
                              .done_ntt(done10_ntt),
                              .f_hat(in_1)
                          );
                          
                          inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_2 (
                              .clk(clk),
                              .rst(rst),
                              .f(mul_add[1]),
                              .start_ntt(start_inverse),
                              .done_ntt(done11_ntt),
                              .f_hat(in_2)
                          );
                          
                          inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_3 (
                              .clk(clk),
                              .rst(rst),
                              .f(mul_add[2]),
                              .start_ntt(start_inverse),
                              .done_ntt(done12_ntt),
                              .f_hat(in_3)
                          );
                           inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_4 (
                                                       .clk(clk),
                                                       .rst(rst),
                                                       .f(mul_add_t[0]),
                                                       .start_ntt(start_inverse),
                                                       .done_ntt(done13_ntt),
                                                       .f_hat(in_4)
                                                   );
                                                   
                        inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_5 (
                                                       .clk(clk),
                                                       .rst(rst),
                                                       .f(mul_add_t[1]),
                                                       .start_ntt(start_inverse),
                                                       .done_ntt(done14_ntt),
                                                       .f_hat(in_5)
                                                   );
                                                   
                        inverse_ntt #(.N(256), .Q(3329), .F(3303)) inverse_6 (
                                                       .clk(clk),
                                                       .rst(rst),
                                                       .f(mul_add_t[2]),
                                                       .start_ntt(start_inverse),
                                                       .done_ntt(done15_ntt),
                                                       .f_hat(in_6)
                                                   );
                           

                      decompress_module decompress_inst0 (
                                            .x(m_dec[0]),
                                            .d(16),
                                            .result(decom_out[0])
                                        );
                                        
                                        decompress_module decompress_inst1 (
                                            .x(m_dec[1]),
                                            .d(16),
                                            .result(decom_out[1])
                                        );
                                        
                                        decompress_module decompress_inst2 (
                                            .x(m_dec[2]),
                                            .d(16),
                                            .result(decom_out[2])
                                        );
                                        
                                        decompress_module decompress_inst3 (
                                            .x(m_dec[3]),
                                            .d(16),
                                            .result(decom_out[3])
                                        );
                                        
                                        decompress_module decompress_inst4 (
                                            .x(m_dec[4]),
                                            .d(16),
                                            .result(decom_out[4])
                                        );
                                        
                                        decompress_module decompress_inst5 (
                                            .x(m_dec[5]),
                                            .d(16),
                                            .result(decom_out[5])
                                        );
                                        
                                        decompress_module decompress_inst6 (
                                            .x(m_dec[6]),
                                            .d(16),
                                            .result(decom_out[6])
                                        );
                                        
                                        decompress_module decompress_inst7 (
                                            .x(m_dec[7]),
                                            .d(16),
                                            .result(decom_out[7])
                                        );
                                        
                                        decompress_module decompress_inst8 (
                                            .x(m_dec[8]),
                                            .d(16),
                                            .result(decom_out[8])
                                        );
                                        
                                        decompress_module decompress_inst9 (
                                            .x(m_dec[9]),
                                            .d(16),
                                            .result(decom_out[9])
                                        );
                                        
                                        decompress_module decompress_inst10 (
                                            .x(m_dec[10]),
                                            .d(16),
                                            .result(decom_out[10])
                                        );
                                        
                                        decompress_module decompress_inst11 (
                                            .x(m_dec[11]),
                                            .d(16),
                                            .result(decom_out[11])
                                        );
                                        
                                        decompress_module decompress_inst12 (
                                            .x(m_dec[12]),
                                            .d(16),
                                            .result(decom_out[12])
                                        );
                                        
                                        decompress_module decompress_inst13 (
                                            .x(m_dec[13]),
                                            .d(16),
                                            .result(decom_out[13])
                                        );
                                        
                                        decompress_module decompress_inst14 (
                                            .x(m_dec[14]),
                                            .d(16),
                                            .result(decom_out[14])
                                        );
                                        
                                        decompress_module decompress_inst15 (
                                            .x(m_dec[15]),
                                            .d(16),
                                            .result(decom_out[15])
                                        );
                                        
                                        decompress_module decompress_inst16 (
                                            .x(m_dec[16]),
                                            .d(16),
                                            .result(decom_out[16])
                                        );
                                        
                                        decompress_module decompress_inst17 (
                                            .x(m_dec[17]),
                                            .d(16),
                                            .result(decom_out[17])
                                        );
                                        
                                        decompress_module decompress_inst18 (
                                            .x(m_dec[18]),
                                            .d(16),
                                            .result(decom_out[18])
                                        );
                                        
                                        decompress_module decompress_inst19 (
                                            .x(m_dec[19]),
                                            .d(16),
                                            .result(decom_out[19])
                                        );
                                        
                                        decompress_module decompress_inst20 (
                                            .x(m_dec[20]),
                                            .d(16),
                                            .result(decom_out[20])
                                        );
                                        
                                        decompress_module decompress_inst21 (
                                            .x(m_dec[21]),
                                            .d(16),
                                            .result(decom_out[21])
                                        );
                                        
                                        decompress_module decompress_inst22 (
                                            .x(m_dec[22]),
                                            .d(16),
                                            .result(decom_out[22])
                                        );
                                        
                                        decompress_module decompress_inst23 (
                                            .x(m_dec[23]),
                                            .d(16),
                                            .result(decom_out[23])
                                        );
                                        
                                        decompress_module decompress_inst24 (
                                            .x(m_dec[24]),
                                            .d(16),
                                            .result(decom_out[24])
                                        );
                                        
                                        decompress_module decompress_inst25 (
                                            .x(m_dec[25]),
                                            .d(16),
                                            .result(decom_out[25])
                                        );
                                        
                                        decompress_module decompress_inst26 (
                                            .x(m_dec[26]),
                                            .d(16),
                                            .result(decom_out[26])
                                        );
                                        
                                        decompress_module decompress_inst27 (
                                            .x(m_dec[27]),
                                            .d(16),
                                            .result(decom_out[27])
                                        );
                                        
                                        decompress_module decompress_inst28 (
                                            .x(m_dec[28]),
                                            .d(16),
                                            .result(decom_out[28])
                                        );
                                        
                                        decompress_module decompress_inst29 (
                                            .x(m_dec[29]),
                                            .d(16),
                                            .result(decom_out[29])
                                        );
                                        
                                        decompress_module decompress_inst30 (
                                            .x(m_dec[30]),
                                            .d(16),
                                            .result(decom_out[30])
                                        );
                                        
                                        decompress_module decompress_inst31 (
                                            .x(m_dec[31]),
                                            .d(16),
                                            .result(decom_out[31])
                                        );
                                        
                                        decompress_module decompress_inst32 (
                                            .x(m_dec[32]),
                                            .d(16),
                                            .result(decom_out[32])
                                        );
                                        
                                        decompress_module decompress_inst33 (
                                            .x(m_dec[33]),
                                            .d(16),
                                            .result(decom_out[33])
                                        );
                                        
                                        decompress_module decompress_inst34 (
                                            .x(m_dec[34]),
                                            .d(16),
                                            .result(decom_out[34])
                                        );
                                        
                                        decompress_module decompress_inst35 (
                                            .x(m_dec[35]),
                                            .d(16),
                                            .result(decom_out[35])
                                        );
                                        
                                        decompress_module decompress_inst36 (
                                            .x(m_dec[36]),
                                            .d(16),
                                            .result(decom_out[36])
                                        );
                                        
                                        decompress_module decompress_inst37 (
                                            .x(m_dec[37]),
                                            .d(16),
                                            .result(decom_out[37])
                                        );
                                        
                                        decompress_module decompress_inst38 (
                                            .x(m_dec[38]),
                                            .d(16),
                                            .result(decom_out[38])
                                        );
                                        
                                        decompress_module decompress_inst39 (
                                            .x(m_dec[39]),
                                            .d(16),
                                            .result(decom_out[39])
                                        );
                                        
                                        decompress_module decompress_inst40 (
                                            .x(m_dec[40]),
                                            .d(16),
                                            .result(decom_out[40])
                                        );
                                        
                                        decompress_module decompress_inst41 (
                                            .x(m_dec[41]),
                                            .d(16),
                                            .result(decom_out[41])
                                        );
                                        
                                        decompress_module decompress_inst42 (
                                            .x(m_dec[42]),
                                            .d(16),
                                            .result(decom_out[42])
                                        );
                                        
                                        decompress_module decompress_inst43 (
                                            .x(m_dec[43]),
                                            .d(16),
                                            .result(decom_out[43])
                                        );
                                        
                                        decompress_module decompress_inst44 (
                                            .x(m_dec[44]),
                                            .d(16),
                                            .result(decom_out[44])
                                        );
                                        
                                        decompress_module decompress_inst45 (
                                            .x(m_dec[45]),
                                            .d(16),
                                            .result(decom_out[45])
                                        );
                                        
                                        decompress_module decompress_inst46 (
                                            .x(m_dec[46]),
                                            .d(16),
                                            .result(decom_out[46])
                                        );
                                        
                                        decompress_module decompress_inst47 (
                                            .x(m_dec[47]),
                                            .d(16),
                                            .result(decom_out[47])
                                        );
                                        
                                        decompress_module decompress_inst48 (
                                            .x(m_dec[48]),
                                            .d(16),
                                            .result(decom_out[48])
                                        );
                                        
                                        decompress_module decompress_inst49 (
                                            .x(m_dec[49]),
                                            .d(16),
                                            .result(decom_out[49])
                                        );
                                        
                                        decompress_module decompress_inst50 (
                                            .x(m_dec[50]),
                                            .d(16),
                                            .result(decom_out[50])
                                        );
                                        
                                        decompress_module decompress_inst51 (
                                            .x(m_dec[51]),
                                            .d(16),
                                            .result(decom_out[51])
                                        );
                                        
                                        decompress_module decompress_inst52 (
                                            .x(m_dec[52]),
                                            .d(16),
                                            .result(decom_out[52])
                                        );
                                        
                                        decompress_module decompress_inst53 (
                                            .x(m_dec[53]),
                                            .d(16),
                                            .result(decom_out[53])
                                        );
                                        
                                        decompress_module decompress_inst54 (
                                            .x(m_dec[54]),
                                            .d(16),
                                            .result(decom_out[54])
                                        );
                                        
                                        decompress_module decompress_inst55 (
                                            .x(m_dec[55]),
                                            .d(16),
                                            .result(decom_out[55])
                                        );
                                        
                                        decompress_module decompress_inst56 (
                                            .x(m_dec[56]),
                                            .d(16),
                                            .result(decom_out[56])
                                        );
                                        
                                        decompress_module decompress_inst57 (
                                            .x(m_dec[57]),
                                            .d(16),
                                            .result(decom_out[57])
                                        );
                                        
                                        decompress_module decompress_inst58 (
                                            .x(m_dec[58]),
                                            .d(16),
                                            .result(decom_out[58])
                                        );
                                        
                                        decompress_module decompress_inst59 (
                                            .x(m_dec[59]),
                                            .d(16),
                                            .result(decom_out[59])
                                        );
                                        
                                        decompress_module decompress_inst60 (
                                            .x(m_dec[60]),
                                            .d(16),
                                            .result(decom_out[60])
                                        );
                                        
                                        decompress_module decompress_inst61 (
                                            .x(m_dec[61]),
                                            .d(16),
                                            .result(decom_out[61])
                                        );
                                        
                                        decompress_module decompress_inst62 (
                                            .x(m_dec[62]),
                                            .d(16),
                                            .result(decom_out[62])
                                        );
                                        
                                        decompress_module decompress_inst63 (
                                            .x(m_dec[63]),
                                            .d(16),
                                            .result(decom_out[63])
                                        );
                                        
                                        decompress_module decompress_inst64 (
                                            .x(m_dec[64]),
                                            .d(16),
                                            .result(decom_out[64])
                                        );
                                        
                                        decompress_module decompress_inst65 (
                                            .x(m_dec[65]),
                                            .d(16),
                                            .result(decom_out[65])
                                        );
                                        
                                        decompress_module decompress_inst66 (
                                            .x(m_dec[66]),
                                            .d(16),
                                            .result(decom_out[66])
                                        );
                                        
                                        decompress_module decompress_inst67 (
                                            .x(m_dec[67]),
                                            .d(16),
                                            .result(decom_out[67])
                                        );
                                        
                                        decompress_module decompress_inst68 (
                                            .x(m_dec[68]),
                                            .d(16),
                                            .result(decom_out[68])
                                        );
                                        
                                        decompress_module decompress_inst69 (
                                            .x(m_dec[69]),
                                            .d(16),
                                            .result(decom_out[69])
                                        );
                                        
                                        decompress_module decompress_inst70 (
                                            .x(m_dec[70]),
                                            .d(16),
                                            .result(decom_out[70])
                                        );
                                        
                                        decompress_module decompress_inst71 (
                                            .x(m_dec[71]),
                                            .d(16),
                                            .result(decom_out[71])
                                        );
                                        
                                        decompress_module decompress_inst72 (
                                            .x(m_dec[72]),
                                            .d(16),
                                            .result(decom_out[72])
                                        );
                                        
                                        decompress_module decompress_inst73 (
                                            .x(m_dec[73]),
                                            .d(16),
                                            .result(decom_out[73])
                                        );
                                        
                                        decompress_module decompress_inst74 (
                                            .x(m_dec[74]),
                                            .d(16),
                                            .result(decom_out[74])
                                        );
                                        
                                        decompress_module decompress_inst75 (
                                            .x(m_dec[75]),
                                            .d(16),
                                            .result(decom_out[75])
                                        );
                                        
                                        decompress_module decompress_inst76 (
                                            .x(m_dec[76]),
                                            .d(16),
                                            .result(decom_out[76])
                                        );
                                        
                                        decompress_module decompress_inst77 (
                                            .x(m_dec[77]),
                                            .d(16),
                                            .result(decom_out[77])
                                        );
                                        
                                        decompress_module decompress_inst78 (
                                            .x(m_dec[78]),
                                            .d(16),
                                            .result(decom_out[78])
                                        );
                                        
                                        decompress_module decompress_inst79 (
                                            .x(m_dec[79]),
                                            .d(16),
                                            .result(decom_out[79])
                                        );
                                        
                                        decompress_module decompress_inst80 (
                                            .x(m_dec[80]),
                                            .d(16),
                                            .result(decom_out[80])
                                        );
                                        
                                        decompress_module decompress_inst81 (
                                            .x(m_dec[81]),
                                            .d(16),
                                            .result(decom_out[81])
                                        );
                                        
                                        decompress_module decompress_inst82 (
                                            .x(m_dec[82]),
                                            .d(16),
                                            .result(decom_out[82])
                                        );
                                        
                                        decompress_module decompress_inst83 (
                                            .x(m_dec[83]),
                                            .d(16),
                                            .result(decom_out[83])
                                        );
                                        
                                        decompress_module decompress_inst84 (
                                            .x(m_dec[84]),
                                            .d(16),
                                            .result(decom_out[84])
                                        );
                                        
                                        decompress_module decompress_inst85 (
                                            .x(m_dec[85]),
                                            .d(16),
                                            .result(decom_out[85])
                                        );
                                        
                                        decompress_module decompress_inst86 (
                                            .x(m_dec[86]),
                                            .d(16),
                                            .result(decom_out[86])
                                        );
                                        
                                        decompress_module decompress_inst87 (
                                            .x(m_dec[87]),
                                            .d(16),
                                            .result(decom_out[87])
                                        );
                                        
                                        decompress_module decompress_inst88 (
                                            .x(m_dec[88]),
                                            .d(16),
                                            .result(decom_out[88])
                                        );
                                        
                                        decompress_module decompress_inst89 (
                                            .x(m_dec[89]),
                                            .d(16),
                                            .result(decom_out[89])
                                        );
                                        
                                        decompress_module decompress_inst90 (
                                            .x(m_dec[90]),
                                            .d(16),
                                            .result(decom_out[90])
                                        );
                                        
                                        decompress_module decompress_inst91 (
                                            .x(m_dec[91]),
                                            .d(16),
                                            .result(decom_out[91])
                                        );
                                        
                                        decompress_module decompress_inst92 (
                                            .x(m_dec[92]),
                                            .d(16),
                                            .result(decom_out[92])
                                        );
                                        
                                        decompress_module decompress_inst93 (
                                            .x(m_dec[93]),
                                            .d(16),
                                            .result(decom_out[93])
                                        );
                                        
                                        decompress_module decompress_inst94 (
                                            .x(m_dec[94]),
                                            .d(16),
                                            .result(decom_out[94])
                                        );
                                        
                                        decompress_module decompress_inst95 (
                                            .x(m_dec[95]),
                                            .d(16),
                                            .result(decom_out[95])
                                        );
                                        
                                        decompress_module decompress_inst96 (
                                            .x(m_dec[96]),
                                            .d(16),
                                            .result(decom_out[96])
                                        );
                                        
                                        decompress_module decompress_inst97 (
                                            .x(m_dec[97]),
                                            .d(16),
                                            .result(decom_out[97])
                                        );
                                        
                                        decompress_module decompress_inst98 (
                                            .x(m_dec[98]),
                                            .d(16),
                                            .result(decom_out[98])
                                        );
                                        
                                        decompress_module decompress_inst99 (
                                            .x(m_dec[99]),
                                            .d(16),
                                            .result(decom_out[99])
                                        );
                                        
                                        decompress_module decompress_inst100 (
                                            .x(m_dec[100]),
                                            .d(16),
                                            .result(decom_out[100])
                                        );
                                        
                                        decompress_module decompress_inst101 (
                                            .x(m_dec[101]),
                                            .d(16),
                                            .result(decom_out[101])
                                        );
                                        
                                        decompress_module decompress_inst102 (
                                            .x(m_dec[102]),
                                            .d(16),
                                            .result(decom_out[102])
                                        );
                                        
                                        decompress_module decompress_inst103 (
                                            .x(m_dec[103]),
                                            .d(16),
                                            .result(decom_out[103])
                                        );
                                        
                                        decompress_module decompress_inst104 (
                                            .x(m_dec[104]),
                                            .d(16),
                                            .result(decom_out[104])
                                        );
                                        
                                        decompress_module decompress_inst105 (
                                            .x(m_dec[105]),
                                            .d(16),
                                            .result(decom_out[105])
                                        );
                                        
                                        decompress_module decompress_inst106 (
                                            .x(m_dec[106]),
                                            .d(16),
                                            .result(decom_out[106])
                                        );
                                        
                                        decompress_module decompress_inst107 (
                                            .x(m_dec[107]),
                                            .d(16),
                                            .result(decom_out[107])
                                        );
                                        
                                        decompress_module decompress_inst108 (
                                            .x(m_dec[108]),
                                            .d(16),
                                            .result(decom_out[108])
                                        );
                                        
                                        decompress_module decompress_inst109 (
                                            .x(m_dec[109]),
                                            .d(16),
                                            .result(decom_out[109])
                                        );
                                        
                                        decompress_module decompress_inst110 (
                                            .x(m_dec[110]),
                                            .d(16),
                                            .result(decom_out[110])
                                        );
                                        
                                        decompress_module decompress_inst111 (
                                            .x(m_dec[111]),
                                            .d(16),
                                            .result(decom_out[111])
                                        );
                                        
                                        decompress_module decompress_inst112 (
                                            .x(m_dec[112]),
                                            .d(16),
                                            .result(decom_out[112])
                                        );
                                        
                                        decompress_module decompress_inst113 (
                                            .x(m_dec[113]),
                                            .d(16),
                                            .result(decom_out[113])
                                        );
                                        
                                        decompress_module decompress_inst114 (
                                            .x(m_dec[114]),
                                            .d(16),
                                            .result(decom_out[114])
                                        );
                                        
                                        decompress_module decompress_inst115 (
                                            .x(m_dec[115]),
                                            .d(16),
                                            .result(decom_out[115])
                                        );
                                        
                                        decompress_module decompress_inst116 (
                                            .x(m_dec[116]),
                                            .d(16),
                                            .result(decom_out[116])
                                        );
                                        
                                        decompress_module decompress_inst117 (
                                            .x(m_dec[117]),
                                            .d(16),
                                            .result(decom_out[117])
                                        );
                                        
                                        decompress_module decompress_inst118 (
                                            .x(m_dec[118]),
                                            .d(16),
                                            .result(decom_out[118])
                                        );
                                        
                                        decompress_module decompress_inst119 (
                                            .x(m_dec[119]),
                                            .d(16),
                                            .result(decom_out[119])
                                        );
                                        
                                        decompress_module decompress_inst120 (
                                            .x(m_dec[120]),
                                            .d(16),
                                            .result(decom_out[120])
                                        );
                                        
                                        decompress_module decompress_inst121 (
                                            .x(m_dec[121]),
                                            .d(16),
                                            .result(decom_out[121])
                                        );
                                        
                                        decompress_module decompress_inst122 (
                                            .x(m_dec[122]),
                                            .d(16),
                                            .result(decom_out[122])
                                        );
                                        
                                        decompress_module decompress_inst123 (
                                            .x(m_dec[123]),
                                            .d(16),
                                            .result(decom_out[123])
                                        );
                                        
                                        decompress_module decompress_inst124 (
                                            .x(m_dec[124]),
                                            .d(16),
                                            .result(decom_out[124])
                                        );
                                        
                                        decompress_module decompress_inst125 (
                                            .x(m_dec[125]),
                                            .d(16),
                                            .result(decom_out[125])
                                        );
                                        
                                        decompress_module decompress_inst126 (
                                            .x(m_dec[126]),
                                            .d(16),
                                            .result(decom_out[126])
                                        );
                                        
                                        decompress_module decompress_inst127 (
                                            .x(m_dec[127]),
                                            .d(16),
                                            .result(decom_out[127])
                                        );
                                        
                                        decompress_module decompress_inst128 (
                                            .x(m_dec[128]),
                                            .d(16),
                                            .result(decom_out[128])
                                        );
                                        
                                        decompress_module decompress_inst129 (
                                            .x(m_dec[129]),
                                            .d(16),
                                            .result(decom_out[129])
                                        );
                                        
                                        decompress_module decompress_inst130 (
                                            .x(m_dec[130]),
                                            .d(16),
                                            .result(decom_out[130])
                                        );
                                        
                                        decompress_module decompress_inst131 (
                                            .x(m_dec[131]),
                                            .d(16),
                                            .result(decom_out[131])
                                        );
                                        
                                        decompress_module decompress_inst132 (
                                            .x(m_dec[132]),
                                            .d(16),
                                            .result(decom_out[132])
                                        );
                                        
                                        decompress_module decompress_inst133 (
                                            .x(m_dec[133]),
                                            .d(16),
                                            .result(decom_out[133])
                                        );
                                        
                                        decompress_module decompress_inst134 (
                                            .x(m_dec[134]),
                                            .d(16),
                                            .result(decom_out[134])
                                        );
                                        
                                        decompress_module decompress_inst135 (
                                            .x(m_dec[135]),
                                            .d(16),
                                            .result(decom_out[135])
                                        );
                                        
                                        decompress_module decompress_inst136 (
                                            .x(m_dec[136]),
                                            .d(16),
                                            .result(decom_out[136])
                                        );
                                        
                                        decompress_module decompress_inst137 (
                                            .x(m_dec[137]),
                                            .d(16),
                                            .result(decom_out[137])
                                        );
                                        
                                        decompress_module decompress_inst138 (
                                            .x(m_dec[138]),
                                            .d(16),
                                            .result(decom_out[138])
                                        );
                                        
                                        decompress_module decompress_inst139 (
                                            .x(m_dec[139]),
                                            .d(16),
                                            .result(decom_out[139])
                                        );
                                        
                                        decompress_module decompress_inst140 (
                                            .x(m_dec[140]),
                                            .d(16),
                                            .result(decom_out[140])
                                        );
                                        
                                        decompress_module decompress_inst141 (
                                            .x(m_dec[141]),
                                            .d(16),
                                            .result(decom_out[141])
                                        );
                                        
                                        decompress_module decompress_inst142 (
                                            .x(m_dec[142]),
                                            .d(16),
                                            .result(decom_out[142])
                                        );
                                        
                                        decompress_module decompress_inst143 (
                                            .x(m_dec[143]),
                                            .d(16),
                                            .result(decom_out[143])
                                        );
                                        
                                        decompress_module decompress_inst144 (
                                            .x(m_dec[144]),
                                            .d(16),
                                            .result(decom_out[144])
                                        );
                                        
                                        decompress_module decompress_inst145 (
                                            .x(m_dec[145]),
                                            .d(16),
                                            .result(decom_out[145])
                                        );
                                        
                                        decompress_module decompress_inst146 (
                                            .x(m_dec[146]),
                                            .d(16),
                                            .result(decom_out[146])
                                        );
                                        
                                        decompress_module decompress_inst147 (
                                            .x(m_dec[147]),
                                            .d(16),
                                            .result(decom_out[147])
                                        );
                                        
                                        decompress_module decompress_inst148 (
                                            .x(m_dec[148]),
                                            .d(16),
                                            .result(decom_out[148])
                                        );
                                        
                                        decompress_module decompress_inst149 (
                                            .x(m_dec[149]),
                                            .d(16),
                                            .result(decom_out[149])
                                        );
                                        
                                        decompress_module decompress_inst150 (
                                            .x(m_dec[150]),
                                            .d(16),
                                            .result(decom_out[150])
                                        );
                                        
                                        decompress_module decompress_inst151 (
                                            .x(m_dec[151]),
                                            .d(16),
                                            .result(decom_out[151])
                                        );
                                        
                                        decompress_module decompress_inst152 (
                                            .x(m_dec[152]),
                                            .d(16),
                                            .result(decom_out[152])
                                        );
                                        
                                        decompress_module decompress_inst153 (
                                            .x(m_dec[153]),
                                            .d(16),
                                            .result(decom_out[153])
                                        );
                                        
                                        decompress_module decompress_inst154 (
                                            .x(m_dec[154]),
                                            .d(16),
                                            .result(decom_out[154])
                                        );
                                        
                                        decompress_module decompress_inst155 (
                                            .x(m_dec[155]),
                                            .d(16),
                                            .result(decom_out[155])
                                        );
                                        
                                        decompress_module decompress_inst156 (
                                            .x(m_dec[156]),
                                            .d(16),
                                            .result(decom_out[156])
                                        );
                                        
                                        decompress_module decompress_inst157 (
                                            .x(m_dec[157]),
                                            .d(16),
                                            .result(decom_out[157])
                                        );
                                        
                                        decompress_module decompress_inst158 (
                                            .x(m_dec[158]),
                                            .d(16),
                                            .result(decom_out[158])
                                        );
                                        
                                        decompress_module decompress_inst159 (
                                            .x(m_dec[159]),
                                            .d(16),
                                            .result(decom_out[159])
                                        );
                                        
                                        decompress_module decompress_inst160 (
                                            .x(m_dec[160]),
                                            .d(16),
                                            .result(decom_out[160])
                                        );
                                        
                                        decompress_module decompress_inst161 (
                                            .x(m_dec[161]),
                                            .d(16),
                                            .result(decom_out[161])
                                        );
                                        
                                        decompress_module decompress_inst162 (
                                            .x(m_dec[162]),
                                            .d(16),
                                            .result(decom_out[162])
                                        );
                                        
                                        decompress_module decompress_inst163 (
                                            .x(m_dec[163]),
                                            .d(16),
                                            .result(decom_out[163])
                                        );
                                        
                                        decompress_module decompress_inst164 (
                                            .x(m_dec[164]),
                                            .d(16),
                                            .result(decom_out[164])
                                        );
                                        
                                        decompress_module decompress_inst165 (
                                            .x(m_dec[165]),
                                            .d(16),
                                            .result(decom_out[165])
                                        );
                                        
                                        decompress_module decompress_inst166 (
                                            .x(m_dec[166]),
                                            .d(16),
                                            .result(decom_out[166])
                                        );
                                        
                                        decompress_module decompress_inst167 (
                                            .x(m_dec[167]),
                                            .d(16),
                                            .result(decom_out[167])
                                        );
                                        
                                        decompress_module decompress_inst168 (
                                            .x(m_dec[168]),
                                            .d(16),
                                            .result(decom_out[168])
                                        );
                                        
                                        decompress_module decompress_inst169 (
                                            .x(m_dec[169]),
                                            .d(16),
                                            .result(decom_out[169])
                                        );
                                        
                                        decompress_module decompress_inst170 (
                                            .x(m_dec[170]),
                                            .d(16),
                                            .result(decom_out[170])
                                        );
                                        
                                        decompress_module decompress_inst171 (
                                            .x(m_dec[171]),
                                            .d(16),
                                            .result(decom_out[171])
                                        );
                                        
                                        decompress_module decompress_inst172 (
                                            .x(m_dec[172]),
                                            .d(16),
                                            .result(decom_out[172])
                                        );
                                        
                                        decompress_module decompress_inst173 (
                                            .x(m_dec[173]),
                                            .d(16),
                                            .result(decom_out[173])
                                        );
                                        
                                        decompress_module decompress_inst174 (
                                            .x(m_dec[174]),
                                            .d(16),
                                            .result(decom_out[174])
                                        );
                                        
                                        decompress_module decompress_inst175 (
                                            .x(m_dec[175]),
                                            .d(16),
                                            .result(decom_out[175])
                                        );
                                        
                                        decompress_module decompress_inst176 (
                                            .x(m_dec[176]),
                                            .d(16),
                                            .result(decom_out[176])
                                        );
                                        
                                        decompress_module decompress_inst177 (
                                            .x(m_dec[177]),
                                            .d(16),
                                            .result(decom_out[177])
                                        );
                                        
                                        decompress_module decompress_inst178 (
                                            .x(m_dec[178]),
                                            .d(16),
                                            .result(decom_out[178])
                                        );
                                        
                                        decompress_module decompress_inst179 (
                                            .x(m_dec[179]),
                                            .d(16),
                                            .result(decom_out[179])
                                        );
                                        
                                        decompress_module decompress_inst180 (
                                            .x(m_dec[180]),
                                            .d(16),
                                            .result(decom_out[180])
                                        );
                                        
                                        decompress_module decompress_inst181 (
                                            .x(m_dec[181]),
                                            .d(16),
                                            .result(decom_out[181])
                                        );
                                        
                                        decompress_module decompress_inst182 (
                                            .x(m_dec[182]),
                                            .d(16),
                                            .result(decom_out[182])
                                        );
                                        
                                        decompress_module decompress_inst183 (
                                            .x(m_dec[183]),
                                            .d(16),
                                            .result(decom_out[183])
                                        );
                                        
                                        decompress_module decompress_inst184 (
                                            .x(m_dec[184]),
                                            .d(16),
                                            .result(decom_out[184])
                                        );
                                        
                                        decompress_module decompress_inst185 (
                                            .x(m_dec[185]),
                                            .d(16),
                                            .result(decom_out[185])
                                        );
                                        
                                        decompress_module decompress_inst186 (
                                            .x(m_dec[186]),
                                            .d(16),
                                            .result(decom_out[186])
                                        );
                                        
                                        decompress_module decompress_inst187 (
                                            .x(m_dec[187]),
                                            .d(16),
                                            .result(decom_out[187])
                                        );
                                        
                                        decompress_module decompress_inst188 (
                                            .x(m_dec[188]),
                                            .d(16),
                                            .result(decom_out[188])
                                        );
                                        
                                        decompress_module decompress_inst189 (
                                            .x(m_dec[189]),
                                            .d(16),
                                            .result(decom_out[189])
                                        );
                                        
                                        decompress_module decompress_inst190 (
                                            .x(m_dec[190]),
                                            .d(16),
                                            .result(decom_out[190])
                                        );
                                        
                                        decompress_module decompress_inst191 (
                                            .x(m_dec[191]),
                                            .d(16),
                                            .result(decom_out[191])
                                        );
                                        
                                        decompress_module decompress_inst192 (
                                            .x(m_dec[192]),
                                            .d(16),
                                            .result(decom_out[192])
                                        );
                                        
                                        decompress_module decompress_inst193 (
                                            .x(m_dec[193]),
                                            .d(16),
                                            .result(decom_out[193])
                                        );
                                        
                                        decompress_module decompress_inst194 (
                                            .x(m_dec[194]),
                                            .d(16),
                                            .result(decom_out[194])
                                        );
                                        
                                        decompress_module decompress_inst195 (
                                            .x(m_dec[195]),
                                            .d(16),
                                            .result(decom_out[195])
                                        );
                                        
                                        decompress_module decompress_inst196 (
                                            .x(m_dec[196]),
                                            .d(16),
                                            .result(decom_out[196])
                                        );
                                        
                                        decompress_module decompress_inst197 (
                                            .x(m_dec[197]),
                                            .d(16),
                                            .result(decom_out[197])
                                        );
                                        
                                        decompress_module decompress_inst198 (
                                            .x(m_dec[198]),
                                            .d(16),
                                            .result(decom_out[198])
                                        );
                                        
                                        decompress_module decompress_inst199 (
                                            .x(m_dec[199]),
                                            .d(16),
                                            .result(decom_out[199])
                                        );
                                        
                                        decompress_module decompress_inst200 (
                                            .x(m_dec[200]),
                                            .d(16),
                                            .result(decom_out[200])
                                        );
                                        
                                        decompress_module decompress_inst201 (
                                            .x(m_dec[201]),
                                            .d(16),
                                            .result(decom_out[201])
                                        );
                                        
                                        decompress_module decompress_inst202 (
                                            .x(m_dec[202]),
                                            .d(16),
                                            .result(decom_out[202])
                                        );
                                        
                                        decompress_module decompress_inst203 (
                                            .x(m_dec[203]),
                                            .d(16),
                                            .result(decom_out[203])
                                        );
                                        
                                        decompress_module decompress_inst204 (
                                            .x(m_dec[204]),
                                            .d(16),
                                            .result(decom_out[204])
                                        );
                                        
                                        decompress_module decompress_inst205 (
                                            .x(m_dec[205]),
                                            .d(16),
                                            .result(decom_out[205])
                                        );
                                        
                                        decompress_module decompress_inst206 (
                                            .x(m_dec[206]),
                                            .d(16),
                                            .result(decom_out[206])
                                        );
                                        
                                        decompress_module decompress_inst207 (
                                            .x(m_dec[207]),
                                            .d(16),
                                            .result(decom_out[207])
                                        );
                                        
                                        decompress_module decompress_inst208 (
                                            .x(m_dec[208]),
                                            .d(16),
                                            .result(decom_out[208])
                                        );
                                        
                                        decompress_module decompress_inst209 (
                                            .x(m_dec[209]),
                                            .d(16),
                                            .result(decom_out[209])
                                        );
                                        
                                        decompress_module decompress_inst210 (
                                            .x(m_dec[210]),
                                            .d(16),
                                            .result(decom_out[210])
                                        );
                                        
                                        decompress_module decompress_inst211 (
                                            .x(m_dec[211]),
                                            .d(16),
                                            .result(decom_out[211])
                                        );
                                        
                                        decompress_module decompress_inst212 (
                                            .x(m_dec[212]),
                                            .d(16),
                                            .result(decom_out[212])
                                        );
                                        
                                        decompress_module decompress_inst213 (
                                            .x(m_dec[213]),
                                            .d(16),
                                            .result(decom_out[213])
                                        );
                                        
                                        decompress_module decompress_inst214 (
                                            .x(m_dec[214]),
                                            .d(16),
                                            .result(decom_out[214])
                                        );
                                        
                                        decompress_module decompress_inst215 (
                                            .x(m_dec[215]),
                                            .d(16),
                                            .result(decom_out[215])
                                        );
                                        
                                        decompress_module decompress_inst216 (
                                            .x(m_dec[216]),
                                            .d(16),
                                            .result(decom_out[216])
                                        );
                                        
                                        decompress_module decompress_inst217 (
                                            .x(m_dec[217]),
                                            .d(16),
                                            .result(decom_out[217])
                                        );
                                        
                                        decompress_module decompress_inst218 (
                                            .x(m_dec[218]),
                                            .d(16),
                                            .result(decom_out[218])
                                        );
                                        
                                        decompress_module decompress_inst219 (
                                            .x(m_dec[219]),
                                            .d(16),
                                            .result(decom_out[219])
                                        );
                                        
                                        decompress_module decompress_inst220 (
                                            .x(m_dec[220]),
                                            .d(16),
                                            .result(decom_out[220])
                                        );
                                        
                                        decompress_module decompress_inst221 (
                                            .x(m_dec[221]),
                                            .d(16),
                                            .result(decom_out[221])
                                        );
                                        
                                        decompress_module decompress_inst222 (
                                            .x(m_dec[222]),
                                            .d(16),
                                            .result(decom_out[222])
                                        );
                                        
                                        decompress_module decompress_inst223 (
                                            .x(m_dec[223]),
                                            .d(16),
                                            .result(decom_out[223])
                                        );
                                        
                                        decompress_module decompress_inst224 (
                                            .x(m_dec[224]),
                                            .d(16),
                                            .result(decom_out[224])
                                        );
                                        
                                        decompress_module decompress_inst225 (
                                            .x(m_dec[225]),
                                            .d(16),
                                            .result(decom_out[225])
                                        );
                                        
                                        decompress_module decompress_inst226 (
                                            .x(m_dec[226]),
                                            .d(16),
                                            .result(decom_out[226])
                                        );
                                        
                                        decompress_module decompress_inst227 (
                                            .x(m_dec[227]),
                                            .d(16),
                                            .result(decom_out[227])
                                        );
                                        
                                        decompress_module decompress_inst228 (
                                            .x(m_dec[228]),
                                            .d(16),
                                            .result(decom_out[228])
                                        );
                                        
                                        decompress_module decompress_inst229 (
                                            .x(m_dec[229]),
                                            .d(16),
                                            .result(decom_out[229])
                                        );
                                        
                                        decompress_module decompress_inst230 (
                                            .x(m_dec[230]),
                                            .d(16),
                                            .result(decom_out[230])
                                        );
                                        
                                        decompress_module decompress_inst231 (
                                            .x(m_dec[231]),
                                            .d(16),
                                            .result(decom_out[231])
                                        );
                                        
                                        decompress_module decompress_inst232 (
                                            .x(m_dec[232]),
                                            .d(16),
                                            .result(decom_out[232])
                                        );
                                        
                                        decompress_module decompress_inst233 (
                                            .x(m_dec[233]),
                                            .d(16),
                                            .result(decom_out[233])
                                        );
                                        
                                        decompress_module decompress_inst234 (
                                            .x(m_dec[234]),
                                            .d(16),
                                            .result(decom_out[234])
                                        );
                                        
                                        decompress_module decompress_inst235 (
                                            .x(m_dec[235]),
                                            .d(16),
                                            .result(decom_out[235])
                                        );
                                        
                                        decompress_module decompress_inst236 (
                                            .x(m_dec[236]),
                                            .d(16),
                                            .result(decom_out[236])
                                        );
                                        
                                        decompress_module decompress_inst237 (
                                            .x(m_dec[237]),
                                            .d(16),
                                            .result(decom_out[237])
                                        );
                                        
                                        decompress_module decompress_inst238 (
                                            .x(m_dec[238]),
                                            .d(16),
                                            .result(decom_out[238])
                                        );
                                        
                                        decompress_module decompress_inst239 (
                                            .x(m_dec[239]),
                                            .d(16),
                                            .result(decom_out[239])
                                        );
                                        
                                        decompress_module decompress_inst240 (
                                            .x(m_dec[240]),
                                            .d(16),
                                            .result(decom_out[240])
                                        );
                                        
                                        decompress_module decompress_inst241 (
                                            .x(m_dec[241]),
                                            .d(16),
                                            .result(decom_out[241])
                                        );
                                        
                                        decompress_module decompress_inst242 (
                                            .x(m_dec[242]),
                                            .d(16),
                                            .result(decom_out[242])
                                        );
                                        
                                        decompress_module decompress_inst243 (
                                            .x(m_dec[243]),
                                            .d(16),
                                            .result(decom_out[243])
                                        );
                                        
                                        decompress_module decompress_inst244 (
                                            .x(m_dec[244]),
                                            .d(16),
                                            .result(decom_out[244])
                                        );
                                        
                                        decompress_module decompress_inst245 (
                                            .x(m_dec[245]),
                                            .d(16),
                                            .result(decom_out[245])
                                        );
                                        
                                        decompress_module decompress_inst246 (
                                            .x(m_dec[246]),
                                            .d(16),
                                            .result(decom_out[246])
                                        );
                                        
                                        decompress_module decompress_inst247 (
                                            .x(m_dec[247]),
                                            .d(16),
                                            .result(decom_out[247])
                                        );
                                        
                                        decompress_module decompress_inst248 (
                                            .x(m_dec[248]),
                                            .d(16),
                                            .result(decom_out[248])
                                        );
                                        
                                        decompress_module decompress_inst249 (
                                            .x(m_dec[249]),
                                            .d(16),
                                            .result(decom_out[249])
                                        );
                                        
                                        decompress_module decompress_inst250 (
                                            .x(m_dec[250]),
                                            .d(16),
                                            .result(decom_out[250])
                                        );
                                        
                                        decompress_module decompress_inst251 (
                                            .x(m_dec[251]),
                                            .d(16),
                                            .result(decom_out[251])
                                        );
                                        
                                        decompress_module decompress_inst252 (
                                            .x(m_dec[252]),
                                            .d(16),
                                            .result(decom_out[252])
                                        );
                                        
                                        decompress_module decompress_inst253 (
                                            .x(m_dec[253]),
                                            .d(16),
                                            .result(decom_out[253])
                                        );
                                        
                                        decompress_module decompress_inst254 (
                                            .x(m_dec[254]),
                                            .d(16),
                                            .result(decom_out[254])
                                        );
                                        
                                        decompress_module decompress_inst255 (
                                            .x(m_dec[255]),
                                            .d(16),
                                            .result(decom_out[255])
                                        );
                                        compress_module compress_0 (
                                            .x(u[0][0]),
                                            .d(10),
                                            .result(com_out[0][0])
                                        );
                                        
                                        compress_module compress_1 (
                                            .x(u[0][1]),
                                            .d(10),
                                            .result(com_out[0][1])
                                        );
                                        
                                        compress_module compress_2 (
                                            .x(u[0][2]),
                                            .d(10),
                                            .result(com_out[0][2])
                                        );
                                        
                                        compress_module compress_3 (
                                            .x(u[0][3]),
                                            .d(10),
                                            .result(com_out[0][3])
                                        );
                                        
                                        compress_module compress_4 (
                                            .x(u[0][4]),
                                            .d(10),
                                            .result(com_out[0][4])
                                        );
                                        
                                        compress_module compress_5 (
                                            .x(u[0][5]),
                                            .d(10),
                                            .result(com_out[0][5])
                                        );
                                        
                                        compress_module compress_6 (
                                            .x(u[0][6]),
                                            .d(10),
                                            .result(com_out[0][6])
                                        );
                                        
                                        compress_module compress_7 (
                                            .x(u[0][7]),
                                            .d(10),
                                            .result(com_out[0][7])
                                        );
                                        
                                        compress_module compress_8 (
                                            .x(u[0][8]),
                                            .d(10),
                                            .result(com_out[0][8])
                                        );
                                        
                                        compress_module compress_9 (
                                            .x(u[0][9]),
                                            .d(10),
                                            .result(com_out[0][9])
                                        );
                                        
                                        compress_module compress_10 (
                                            .x(u[0][10]),
                                            .d(10),
                                            .result(com_out[0][10])
                                        );
                                        
                                        compress_module compress_11 (
                                            .x(u[0][11]),
                                            .d(10),
                                            .result(com_out[0][11])
                                        );
                                        
                                        compress_module compress_12 (
                                            .x(u[0][12]),
                                            .d(10),
                                            .result(com_out[0][12])
                                        );
                                        
                                        compress_module compress_13 (
                                            .x(u[0][13]),
                                            .d(10),
                                            .result(com_out[0][13])
                                        );
                                        
                                        compress_module compress_14 (
                                            .x(u[0][14]),
                                            .d(10),
                                            .result(com_out[0][14])
                                        );
                                        
                                        compress_module compress_15 (
                                            .x(u[0][15]),
                                            .d(10),
                                            .result(com_out[0][15])
                                        );
                                        
                                        compress_module compress_16 (
                                            .x(u[0][16]),
                                            .d(10),
                                            .result(com_out[0][16])
                                        );
                                        
                                        compress_module compress_17 (
                                            .x(u[0][17]),
                                            .d(10),
                                            .result(com_out[0][17])
                                        );
                                        
                                        compress_module compress_18 (
                                            .x(u[0][18]),
                                            .d(10),
                                            .result(com_out[0][18])
                                        );
                                        
                                        compress_module compress_19 (
                                            .x(u[0][19]),
                                            .d(10),
                                            .result(com_out[0][19])
                                        );
                                        
                                        compress_module compress_20 (
                                            .x(u[0][20]),
                                            .d(10),
                                            .result(com_out[0][20])
                                        );
                                        
                                        compress_module compress_21 (
                                            .x(u[0][21]),
                                            .d(10),
                                            .result(com_out[0][21])
                                        );
                                        
                                        compress_module compress_22 (
                                            .x(u[0][22]),
                                            .d(10),
                                            .result(com_out[0][22])
                                        );
                                        
                                        compress_module compress_23 (
                                            .x(u[0][23]),
                                            .d(10),
                                            .result(com_out[0][23])
                                        );
                                        
                                        compress_module compress_24 (
                                            .x(u[0][24]),
                                            .d(10),
                                            .result(com_out[0][24])
                                        );
                                        
                                        compress_module compress_25 (
                                            .x(u[0][25]),
                                            .d(10),
                                            .result(com_out[0][25])
                                        );
                                        
                                        compress_module compress_26 (
                                            .x(u[0][26]),
                                            .d(10),
                                            .result(com_out[0][26])
                                        );
                                        
                                        compress_module compress_27 (
                                            .x(u[0][27]),
                                            .d(10),
                                            .result(com_out[0][27])
                                        );
                                        
                                        compress_module compress_28 (
                                            .x(u[0][28]),
                                            .d(10),
                                            .result(com_out[0][28])
                                        );
                                        
                                        compress_module compress_29 (
                                            .x(u[0][29]),
                                            .d(10),
                                            .result(com_out[0][29])
                                        );
                                        
                                        compress_module compress_30 (
                                            .x(u[0][30]),
                                            .d(10),
                                            .result(com_out[0][30])
                                        );
                                        
                                        compress_module compress_31 (
                                            .x(u[0][31]),
                                            .d(10),
                                            .result(com_out[0][31])
                                        );
                                        
                                        compress_module compress_32 (
                                            .x(u[0][32]),
                                            .d(10),
                                            .result(com_out[0][32])
                                        );
                                        
                                        compress_module compress_33 (
                                            .x(u[0][33]),
                                            .d(10),
                                            .result(com_out[0][33])
                                        );
                                        
                                        compress_module compress_34 (
                                            .x(u[0][34]),
                                            .d(10),
                                            .result(com_out[0][34])
                                        );
                                        
                                        compress_module compress_35 (
                                            .x(u[0][35]),
                                            .d(10),
                                            .result(com_out[0][35])
                                        );
                                        
                                        compress_module compress_36 (
                                            .x(u[0][36]),
                                            .d(10),
                                            .result(com_out[0][36])
                                        );
                                        
                                        compress_module compress_37 (
                                            .x(u[0][37]),
                                            .d(10),
                                            .result(com_out[0][37])
                                        );
                                        
                                        compress_module compress_38 (
                                            .x(u[0][38]),
                                            .d(10),
                                            .result(com_out[0][38])
                                        );
                                        
                                        compress_module compress_39 (
                                            .x(u[0][39]),
                                            .d(10),
                                            .result(com_out[0][39])
                                        );
                                        
                                        compress_module compress_40 (
                                            .x(u[0][40]),
                                            .d(10),
                                            .result(com_out[0][40])
                                        );
                                        
                                        compress_module compress_41 (
                                            .x(u[0][41]),
                                            .d(10),
                                            .result(com_out[0][41])
                                        );
                                        
                                        compress_module compress_42 (
                                            .x(u[0][42]),
                                            .d(10),
                                            .result(com_out[0][42])
                                        );
                                        
                                        compress_module compress_43 (
                                            .x(u[0][43]),
                                            .d(10),
                                            .result(com_out[0][43])
                                        );
                                        
                                        compress_module compress_44 (
                                            .x(u[0][44]),
                                            .d(10),
                                            .result(com_out[0][44])
                                        );
                                        
                                        compress_module compress_45 (
                                            .x(u[0][45]),
                                            .d(10),
                                            .result(com_out[0][45])
                                        );
                                        
                                        compress_module compress_46 (
                                            .x(u[0][46]),
                                            .d(10),
                                            .result(com_out[0][46])
                                        );
                                        
                                        compress_module compress_47 (
                                            .x(u[0][47]),
                                            .d(10),
                                            .result(com_out[0][47])
                                        );
                                        
                                        compress_module compress_48 (
                                            .x(u[0][48]),
                                            .d(10),
                                            .result(com_out[0][48])
                                        );
                                        
                                        compress_module compress_49 (
                                            .x(u[0][49]),
                                            .d(10),
                                            .result(com_out[0][49])
                                        );
                                        
                                        compress_module compress_50 (
                                            .x(u[0][50]),
                                            .d(10),
                                            .result(com_out[0][50])
                                        );
                                        
                                        compress_module compress_51 (
                                            .x(u[0][51]),
                                            .d(10),
                                            .result(com_out[0][51])
                                        );
                                        
                                        compress_module compress_52 (
                                            .x(u[0][52]),
                                            .d(10),
                                            .result(com_out[0][52])
                                        );
                                        
                                        compress_module compress_53 (
                                            .x(u[0][53]),
                                            .d(10),
                                            .result(com_out[0][53])
                                        );
                                        
                                        compress_module compress_54 (
                                            .x(u[0][54]),
                                            .d(10),
                                            .result(com_out[0][54])
                                        );
                                        
                                        compress_module compress_55 (
                                            .x(u[0][55]),
                                            .d(10),
                                            .result(com_out[0][55])
                                        );
                                        
                                        compress_module compress_56 (
                                            .x(u[0][56]),
                                            .d(10),
                                            .result(com_out[0][56])
                                        );
                                        
                                        compress_module compress_57 (
                                            .x(u[0][57]),
                                            .d(10),
                                            .result(com_out[0][57])
                                        );
                                        
                                        compress_module compress_58 (
                                            .x(u[0][58]),
                                            .d(10),
                                            .result(com_out[0][58])
                                        );
                                        
                                        compress_module compress_59 (
                                            .x(u[0][59]),
                                            .d(10),
                                            .result(com_out[0][59])
                                        );
                                        
                                        compress_module compress_60 (
                                            .x(u[0][60]),
                                            .d(10),
                                            .result(com_out[0][60])
                                        );
                                        
                                        compress_module compress_61 (
                                            .x(u[0][61]),
                                            .d(10),
                                            .result(com_out[0][61])
                                        );
                                        
                                        compress_module compress_62 (
                                            .x(u[0][62]),
                                            .d(10),
                                            .result(com_out[0][62])
                                        );
                                        
                                        compress_module compress_63 (
                                            .x(u[0][63]),
                                            .d(10),
                                            .result(com_out[0][63])
                                        );
                                        
                                        compress_module compress_64 (
                                            .x(u[0][64]),
                                            .d(10),
                                            .result(com_out[0][64])
                                        );
                                        
                                        compress_module compress_65 (
                                            .x(u[0][65]),
                                            .d(10),
                                            .result(com_out[0][65])
                                        );
                                        
                                        compress_module compress_66 (
                                            .x(u[0][66]),
                                            .d(10),
                                            .result(com_out[0][66])
                                        );
                                        
                                        compress_module compress_67 (
                                            .x(u[0][67]),
                                            .d(10),
                                            .result(com_out[0][67])
                                        );
                                        
                                        compress_module compress_68 (
                                            .x(u[0][68]),
                                            .d(10),
                                            .result(com_out[0][68])
                                        );
                                        
                                        compress_module compress_69 (
                                            .x(u[0][69]),
                                            .d(10),
                                            .result(com_out[0][69])
                                        );
                                        
                                        compress_module compress_70 (
                                            .x(u[0][70]),
                                            .d(10),
                                            .result(com_out[0][70])
                                        );
                                        
                                        compress_module compress_71 (
                                            .x(u[0][71]),
                                            .d(10),
                                            .result(com_out[0][71])
                                        );
                                        
                                        compress_module compress_72 (
                                            .x(u[0][72]),
                                            .d(10),
                                            .result(com_out[0][72])
                                        );
                                        
                                        compress_module compress_73 (
                                            .x(u[0][73]),
                                            .d(10),
                                            .result(com_out[0][73])
                                        );
                                        
                                        compress_module compress_74 (
                                            .x(u[0][74]),
                                            .d(10),
                                            .result(com_out[0][74])
                                        );
                                        
                                        compress_module compress_75 (
                                            .x(u[0][75]),
                                            .d(10),
                                            .result(com_out[0][75])
                                        );
                                        
                                        compress_module compress_76 (
                                            .x(u[0][76]),
                                            .d(10),
                                            .result(com_out[0][76])
                                        );
                                        
                                        compress_module compress_77 (
                                            .x(u[0][77]),
                                            .d(10),
                                            .result(com_out[0][77])
                                        );
                                        
                                        compress_module compress_78 (
                                            .x(u[0][78]),
                                            .d(10),
                                            .result(com_out[0][78])
                                        );
                                        
                                        compress_module compress_79 (
                                            .x(u[0][79]),
                                            .d(10),
                                            .result(com_out[0][79])
                                        );
                                        
                                        compress_module compress_80 (
                                            .x(u[0][80]),
                                            .d(10),
                                            .result(com_out[0][80])
                                        );
                                        
                                        compress_module compress_81 (
                                            .x(u[0][81]),
                                            .d(10),
                                            .result(com_out[0][81])
                                        );
                                        
                                        compress_module compress_82 (
                                            .x(u[0][82]),
                                            .d(10),
                                            .result(com_out[0][82])
                                        );
                                        
                                        compress_module compress_83 (
                                            .x(u[0][83]),
                                            .d(10),
                                            .result(com_out[0][83])
                                        );
                                        
                                        compress_module compress_84 (
                                            .x(u[0][84]),
                                            .d(10),
                                            .result(com_out[0][84])
                                        );
                                        
                                        compress_module compress_85 (
                                            .x(u[0][85]),
                                            .d(10),
                                            .result(com_out[0][85])
                                        );
                                        
                                        compress_module compress_86 (
                                            .x(u[0][86]),
                                            .d(10),
                                            .result(com_out[0][86])
                                        );
                                        
                                        compress_module compress_87 (
                                            .x(u[0][87]),
                                            .d(10),
                                            .result(com_out[0][87])
                                        );
                                        
                                        compress_module compress_88 (
                                            .x(u[0][88]),
                                            .d(10),
                                            .result(com_out[0][88])
                                        );
                                        
                                        compress_module compress_89 (
                                            .x(u[0][89]),
                                            .d(10),
                                            .result(com_out[0][89])
                                        );
                                        
                                        compress_module compress_90 (
                                            .x(u[0][90]),
                                            .d(10),
                                            .result(com_out[0][90])
                                        );
                                        
                                        compress_module compress_91 (
                                            .x(u[0][91]),
                                            .d(10),
                                            .result(com_out[0][91])
                                        );
                                        
                                        compress_module compress_92 (
                                            .x(u[0][92]),
                                            .d(10),
                                            .result(com_out[0][92])
                                        );
                                        
                                        compress_module compress_93 (
                                            .x(u[0][93]),
                                            .d(10),
                                            .result(com_out[0][93])
                                        );
                                        
                                        compress_module compress_94 (
                                            .x(u[0][94]),
                                            .d(10),
                                            .result(com_out[0][94])
                                        );
                                        
                                        compress_module compress_95 (
                                            .x(u[0][95]),
                                            .d(10),
                                            .result(com_out[0][95])
                                        );
                                        
                                        compress_module compress_96 (
                                            .x(u[0][96]),
                                            .d(10),
                                            .result(com_out[0][96])
                                        );
                                        
                                        compress_module compress_97 (
                                            .x(u[0][97]),
                                            .d(10),
                                            .result(com_out[0][97])
                                        );
                                        
                                        compress_module compress_98 (
                                            .x(u[0][98]),
                                            .d(10),
                                            .result(com_out[0][98])
                                        );
                                        
                                        compress_module compress_99 (
                                            .x(u[0][99]),
                                            .d(10),
                                            .result(com_out[0][99])
                                        );
                                        
                                        compress_module compress_100 (
                                            .x(u[0][100]),
                                            .d(10),
                                            .result(com_out[0][100])
                                        );
                                        
                                        compress_module compress_101 (
                                            .x(u[0][101]),
                                            .d(10),
                                            .result(com_out[0][101])
                                        );
                                        
                                        compress_module compress_102 (
                                            .x(u[0][102]),
                                            .d(10),
                                            .result(com_out[0][102])
                                        );
                                        
                                        compress_module compress_103 (
                                            .x(u[0][103]),
                                            .d(10),
                                            .result(com_out[0][103])
                                        );
                                        
                                        compress_module compress_104 (
                                            .x(u[0][104]),
                                            .d(10),
                                            .result(com_out[0][104])
                                        );
                                        
                                        compress_module compress_105 (
                                            .x(u[0][105]),
                                            .d(10),
                                            .result(com_out[0][105])
                                        );
                                        
                                        compress_module compress_106 (
                                            .x(u[0][106]),
                                            .d(10),
                                            .result(com_out[0][106])
                                        );
                                        
                                        compress_module compress_107 (
                                            .x(u[0][107]),
                                            .d(10),
                                            .result(com_out[0][107])
                                        );
                                        
                                        compress_module compress_108 (
                                            .x(u[0][108]),
                                            .d(10),
                                            .result(com_out[0][108])
                                        );
                                        
                                        compress_module compress_109 (
                                            .x(u[0][109]),
                                            .d(10),
                                            .result(com_out[0][109])
                                        );
                                        
                                        compress_module compress_110 (
                                            .x(u[0][110]),
                                            .d(10),
                                            .result(com_out[0][110])
                                        );
                                        
                                        compress_module compress_111 (
                                            .x(u[0][111]),
                                            .d(10),
                                            .result(com_out[0][111])
                                        );
                                        
                                        compress_module compress_112 (
                                            .x(u[0][112]),
                                            .d(10),
                                            .result(com_out[0][112])
                                        );
                                        
                                        compress_module compress_113 (
                                            .x(u[0][113]),
                                            .d(10),
                                            .result(com_out[0][113])
                                        );
                                        
                                        compress_module compress_114 (
                                            .x(u[0][114]),
                                            .d(10),
                                            .result(com_out[0][114])
                                        );
                                        
                                        compress_module compress_115 (
                                            .x(u[0][115]),
                                            .d(10),
                                            .result(com_out[0][115])
                                        );
                                        
                                        compress_module compress_116 (
                                            .x(u[0][116]),
                                            .d(10),
                                            .result(com_out[0][116])
                                        );
                                        
                                        compress_module compress_117 (
                                            .x(u[0][117]),
                                            .d(10),
                                            .result(com_out[0][117])
                                        );
                                        
                                        compress_module compress_118 (
                                            .x(u[0][118]),
                                            .d(10),
                                            .result(com_out[0][118])
                                        );
                                        
                                        compress_module compress_119 (
                                            .x(u[0][119]),
                                            .d(10),
                                            .result(com_out[0][119])
                                        );
                                        
                                        compress_module compress_120 (
                                            .x(u[0][120]),
                                            .d(10),
                                            .result(com_out[0][120])
                                        );
                                        
                                        compress_module compress_121 (
                                            .x(u[0][121]),
                                            .d(10),
                                            .result(com_out[0][121])
                                        );
                                        
                                        compress_module compress_122 (
                                            .x(u[0][122]),
                                            .d(10),
                                            .result(com_out[0][122])
                                        );
                                        
                                        compress_module compress_123 (
                                            .x(u[0][123]),
                                            .d(10),
                                            .result(com_out[0][123])
                                        );
                                        
                                        compress_module compress_124 (
                                            .x(u[0][124]),
                                            .d(10),
                                            .result(com_out[0][124])
                                        );
                                        
                                        compress_module compress_125 (
                                            .x(u[0][125]),
                                            .d(10),
                                            .result(com_out[0][125])
                                        );
                                        
                                        compress_module compress_126 (
                                            .x(u[0][126]),
                                            .d(10),
                                            .result(com_out[0][126])
                                        );
                                        
                                        compress_module compress_127 (
                                            .x(u[0][127]),
                                            .d(10),
                                            .result(com_out[0][127])
                                        );
                                        
                                        compress_module compress_128 (
                                            .x(u[0][128]),
                                            .d(10),
                                            .result(com_out[0][128])
                                        );
                                        
                                        compress_module compress_129 (
                                            .x(u[0][129]),
                                            .d(10),
                                            .result(com_out[0][129])
                                        );
                                        
                                        compress_module compress_130 (
                                            .x(u[0][130]),
                                            .d(10),
                                            .result(com_out[0][130])
                                        );
                                        
                                        compress_module compress_131 (
                                            .x(u[0][131]),
                                            .d(10),
                                            .result(com_out[0][131])
                                        );
                                        
                                        compress_module compress_132 (
                                            .x(u[0][132]),
                                            .d(10),
                                            .result(com_out[0][132])
                                        );
                                        
                                        compress_module compress_133 (
                                            .x(u[0][133]),
                                            .d(10),
                                            .result(com_out[0][133])
                                        );
                                        
                                        compress_module compress_134 (
                                            .x(u[0][134]),
                                            .d(10),
                                            .result(com_out[0][134])
                                        );
                                        
                                        compress_module compress_135 (
                                            .x(u[0][135]),
                                            .d(10),
                                            .result(com_out[0][135])
                                        );
                                        
                                        compress_module compress_136 (
                                            .x(u[0][136]),
                                            .d(10),
                                            .result(com_out[0][136])
                                        );
                                        
                                        compress_module compress_137 (
                                            .x(u[0][137]),
                                            .d(10),
                                            .result(com_out[0][137])
                                        );
                                        
                                        compress_module compress_138 (
                                            .x(u[0][138]),
                                            .d(10),
                                            .result(com_out[0][138])
                                        );
                                        
                                        compress_module compress_139 (
                                            .x(u[0][139]),
                                            .d(10),
                                            .result(com_out[0][139])
                                        );
                                        
                                        compress_module compress_140 (
                                            .x(u[0][140]),
                                            .d(10),
                                            .result(com_out[0][140])
                                        );
                                        
                                        compress_module compress_141 (
                                            .x(u[0][141]),
                                            .d(10),
                                            .result(com_out[0][141])
                                        );
                                        
                                        compress_module compress_142 (
                                            .x(u[0][142]),
                                            .d(10),
                                            .result(com_out[0][142])
                                        );
                                        
                                        compress_module compress_143 (
                                            .x(u[0][143]),
                                            .d(10),
                                            .result(com_out[0][143])
                                        );
                                        
                                        compress_module compress_144 (
                                            .x(u[0][144]),
                                            .d(10),
                                            .result(com_out[0][144])
                                        );
                                        
                                        compress_module compress_145 (
                                            .x(u[0][145]),
                                            .d(10),
                                            .result(com_out[0][145])
                                        );
                                        
                                        compress_module compress_146 (
                                            .x(u[0][146]),
                                            .d(10),
                                            .result(com_out[0][146])
                                        );
                                        
                                        compress_module compress_147 (
                                            .x(u[0][147]),
                                            .d(10),
                                            .result(com_out[0][147])
                                        );
                                        
                                        compress_module compress_148 (
                                            .x(u[0][148]),
                                            .d(10),
                                            .result(com_out[0][148])
                                        );
                                        
                                        compress_module compress_149 (
                                            .x(u[0][149]),
                                            .d(10),
                                            .result(com_out[0][149])
                                        );
                                        
                                        compress_module compress_150 (
                                            .x(u[0][150]),
                                            .d(10),
                                            .result(com_out[0][150])
                                        );
                                        
                                        compress_module compress_151 (
                                            .x(u[0][151]),
                                            .d(10),
                                            .result(com_out[0][151])
                                        );
                                        
                                        compress_module compress_152 (
                                            .x(u[0][152]),
                                            .d(10),
                                            .result(com_out[0][152])
                                        );
                                        
                                        compress_module compress_153 (
                                            .x(u[0][153]),
                                            .d(10),
                                            .result(com_out[0][153])
                                        );
                                        
                                        compress_module compress_154 (
                                            .x(u[0][154]),
                                            .d(10),
                                            .result(com_out[0][154])
                                        );
                                        
                                        compress_module compress_155 (
                                            .x(u[0][155]),
                                            .d(10),
                                            .result(com_out[0][155])
                                        );
                                        
                                        compress_module compress_156 (
                                            .x(u[0][156]),
                                            .d(10),
                                            .result(com_out[0][156])
                                        );
                                        
                                        compress_module compress_157 (
                                            .x(u[0][157]),
                                            .d(10),
                                            .result(com_out[0][157])
                                        );
                                        
                                        compress_module compress_158 (
                                            .x(u[0][158]),
                                            .d(10),
                                            .result(com_out[0][158])
                                        );
                                        
                                        compress_module compress_159 (
                                            .x(u[0][159]),
                                            .d(10),
                                            .result(com_out[0][159])
                                        );
                                        
                                        compress_module compress_160 (
                                            .x(u[0][160]),
                                            .d(10),
                                            .result(com_out[0][160])
                                        );
                                        
                                        compress_module compress_161 (
                                            .x(u[0][161]),
                                            .d(10),
                                            .result(com_out[0][161])
                                        );
                                        
                                        compress_module compress_162 (
                                            .x(u[0][162]),
                                            .d(10),
                                            .result(com_out[0][162])
                                        );
                                        
                                        compress_module compress_163 (
                                            .x(u[0][163]),
                                            .d(10),
                                            .result(com_out[0][163])
                                        );
                                        
                                        compress_module compress_164 (
                                            .x(u[0][164]),
                                            .d(10),
                                            .result(com_out[0][164])
                                        );
                                        
                                        compress_module compress_165 (
                                            .x(u[0][165]),
                                            .d(10),
                                            .result(com_out[0][165])
                                        );
                                        
                                        compress_module compress_166 (
                                            .x(u[0][166]),
                                            .d(10),
                                            .result(com_out[0][166])
                                        );
                                        
                                        compress_module compress_167 (
                                            .x(u[0][167]),
                                            .d(10),
                                            .result(com_out[0][167])
                                        );
                                        
                                        compress_module compress_168 (
                                            .x(u[0][168]),
                                            .d(10),
                                            .result(com_out[0][168])
                                        );
                                        
                                        compress_module compress_169 (
                                            .x(u[0][169]),
                                            .d(10),
                                            .result(com_out[0][169])
                                        );
                                        
                                        compress_module compress_170 (
                                            .x(u[0][170]),
                                            .d(10),
                                            .result(com_out[0][170])
                                        );
                                        
                                        compress_module compress_171 (
                                            .x(u[0][171]),
                                            .d(10),
                                            .result(com_out[0][171])
                                        );
                                        
                                        compress_module compress_172 (
                                            .x(u[0][172]),
                                            .d(10),
                                            .result(com_out[0][172])
                                        );
                                        
                                        compress_module compress_173 (
                                            .x(u[0][173]),
                                            .d(10),
                                            .result(com_out[0][173])
                                        );
                                        
                                        compress_module compress_174 (
                                            .x(u[0][174]),
                                            .d(10),
                                            .result(com_out[0][174])
                                        );
                                        
                                        compress_module compress_175 (
                                            .x(u[0][175]),
                                            .d(10),
                                            .result(com_out[0][175])
                                        );
                                        
                                        compress_module compress_176 (
                                            .x(u[0][176]),
                                            .d(10),
                                            .result(com_out[0][176])
                                        );
                                        
                                        compress_module compress_177 (
                                            .x(u[0][177]),
                                            .d(10),
                                            .result(com_out[0][177])
                                        );
                                        
                                        compress_module compress_178 (
                                            .x(u[0][178]),
                                            .d(10),
                                            .result(com_out[0][178])
                                        );
                                        
                                        compress_module compress_179 (
                                            .x(u[0][179]),
                                            .d(10),
                                            .result(com_out[0][179])
                                        );
                                        
                                        compress_module compress_180 (
                                            .x(u[0][180]),
                                            .d(10),
                                            .result(com_out[0][180])
                                        );
                                        
                                        compress_module compress_181 (
                                            .x(u[0][181]),
                                            .d(10),
                                            .result(com_out[0][181])
                                        );
                                        
                                        compress_module compress_182 (
                                            .x(u[0][182]),
                                            .d(10),
                                            .result(com_out[0][182])
                                        );
                                        
                                        compress_module compress_183 (
                                            .x(u[0][183]),
                                            .d(10),
                                            .result(com_out[0][183])
                                        );
                                        
                                        compress_module compress_184 (
                                            .x(u[0][184]),
                                            .d(10),
                                            .result(com_out[0][184])
                                        );
                                        
                                        compress_module compress_185 (
                                            .x(u[0][185]),
                                            .d(10),
                                            .result(com_out[0][185])
                                        );
                                        
                                        compress_module compress_186 (
                                            .x(u[0][186]),
                                            .d(10),
                                            .result(com_out[0][186])
                                        );
                                        
                                        compress_module compress_187 (
                                            .x(u[0][187]),
                                            .d(10),
                                            .result(com_out[0][187])
                                        );
                                        
                                        compress_module compress_188 (
                                            .x(u[0][188]),
                                            .d(10),
                                            .result(com_out[0][188])
                                        );
                                        
                                        compress_module compress_189 (
                                            .x(u[0][189]),
                                            .d(10),
                                            .result(com_out[0][189])
                                        );
                                        
                                        compress_module compress_190 (
                                            .x(u[0][190]),
                                            .d(10),
                                            .result(com_out[0][190])
                                        );
                                        
                                        compress_module compress_191 (
                                            .x(u[0][191]),
                                            .d(10),
                                            .result(com_out[0][191])
                                        );
                                        
                                        compress_module compress_192 (
                                            .x(u[0][192]),
                                            .d(10),
                                            .result(com_out[0][192])
                                        );
                                        
                                        compress_module compress_193 (
                                            .x(u[0][193]),
                                            .d(10),
                                            .result(com_out[0][193])
                                        );
                                        
                                        compress_module compress_194 (
                                            .x(u[0][194]),
                                            .d(10),
                                            .result(com_out[0][194])
                                        );
                                        
                                        compress_module compress_195 (
                                            .x(u[0][195]),
                                            .d(10),
                                            .result(com_out[0][195])
                                        );
                                        
                                        compress_module compress_196 (
                                            .x(u[0][196]),
                                            .d(10),
                                            .result(com_out[0][196])
                                        );
                                        
                                        compress_module compress_197 (
                                            .x(u[0][197]),
                                            .d(10),
                                            .result(com_out[0][197])
                                        );
                                        
                                        compress_module compress_198 (
                                            .x(u[0][198]),
                                            .d(10),
                                            .result(com_out[0][198])
                                        );
                                        
                                        compress_module compress_199 (
                                            .x(u[0][199]),
                                            .d(10),
                                            .result(com_out[0][199])
                                        );
                                        
                                        compress_module compress_200 (
                                            .x(u[0][200]),
                                            .d(10),
                                            .result(com_out[0][200])
                                        );
                                        
                                        compress_module compress_201 (
                                            .x(u[0][201]),
                                            .d(10),
                                            .result(com_out[0][201])
                                        );
                                        
                                        compress_module compress_202 (
                                            .x(u[0][202]),
                                            .d(10),
                                            .result(com_out[0][202])
                                        );
                                        
                                        compress_module compress_203 (
                                            .x(u[0][203]),
                                            .d(10),
                                            .result(com_out[0][203])
                                        );
                                        
                                        compress_module compress_204 (
                                            .x(u[0][204]),
                                            .d(10),
                                            .result(com_out[0][204])
                                        );
                                        
                                        compress_module compress_205 (
                                            .x(u[0][205]),
                                            .d(10),
                                            .result(com_out[0][205])
                                        );
                                        
                                        compress_module compress_206 (
                                            .x(u[0][206]),
                                            .d(10),
                                            .result(com_out[0][206])
                                        );
                                        
                                        compress_module compress_207 (
                                            .x(u[0][207]),
                                            .d(10),
                                            .result(com_out[0][207])
                                        );
                                        
                                        compress_module compress_208 (
                                            .x(u[0][208]),
                                            .d(10),
                                            .result(com_out[0][208])
                                        );
                                        
                                        compress_module compress_209 (
                                            .x(u[0][209]),
                                            .d(10),
                                            .result(com_out[0][209])
                                        );
                                        
                                        compress_module compress_210 (
                                            .x(u[0][210]),
                                            .d(10),
                                            .result(com_out[0][210])
                                        );
                                        
                                        compress_module compress_211 (
                                            .x(u[0][211]),
                                            .d(10),
                                            .result(com_out[0][211])
                                        );
                                        
                                        compress_module compress_212 (
                                            .x(u[0][212]),
                                            .d(10),
                                            .result(com_out[0][212])
                                        );
                                        
                                        compress_module compress_213 (
                                            .x(u[0][213]),
                                            .d(10),
                                            .result(com_out[0][213])
                                        );
                                        
                                        compress_module compress_214 (
                                            .x(u[0][214]),
                                            .d(10),
                                            .result(com_out[0][214])
                                        );
                                        
                                        compress_module compress_215 (
                                            .x(u[0][215]),
                                            .d(10),
                                            .result(com_out[0][215])
                                        );
                                        
                                        compress_module compress_216 (
                                            .x(u[0][216]),
                                            .d(10),
                                            .result(com_out[0][216])
                                        );
                                        
                                        compress_module compress_217 (
                                            .x(u[0][217]),
                                            .d(10),
                                            .result(com_out[0][217])
                                        );
                                        
                                        compress_module compress_218 (
                                            .x(u[0][218]),
                                            .d(10),
                                            .result(com_out[0][218])
                                        );
                                        
                                        compress_module compress_219 (
                                            .x(u[0][219]),
                                            .d(10),
                                            .result(com_out[0][219])
                                        );
                                        
                                        compress_module compress_220 (
                                            .x(u[0][220]),
                                            .d(10),
                                            .result(com_out[0][220])
                                        );
                                        
                                        compress_module compress_221 (
                                            .x(u[0][221]),
                                            .d(10),
                                            .result(com_out[0][221])
                                        );
                                        
                                        compress_module compress_222 (
                                            .x(u[0][222]),
                                            .d(10),
                                            .result(com_out[0][222])
                                        );
                                        
                                        compress_module compress_223 (
                                            .x(u[0][223]),
                                            .d(10),
                                            .result(com_out[0][223])
                                        );
                                        
                                        compress_module compress_224 (
                                            .x(u[0][224]),
                                            .d(10),
                                            .result(com_out[0][224])
                                        );
                                        
                                        compress_module compress_225 (
                                            .x(u[0][225]),
                                            .d(10),
                                            .result(com_out[0][225])
                                        );
                                        
                                        compress_module compress_226 (
                                            .x(u[0][226]),
                                            .d(10),
                                            .result(com_out[0][226])
                                        );
                                        
                                        compress_module compress_227 (
                                            .x(u[0][227]),
                                            .d(10),
                                            .result(com_out[0][227])
                                        );
                                        
                                        compress_module compress_228 (
                                            .x(u[0][228]),
                                            .d(10),
                                            .result(com_out[0][228])
                                        );
                                        
                                        compress_module compress_229 (
                                            .x(u[0][229]),
                                            .d(10),
                                            .result(com_out[0][229])
                                        );
                                        
                                        compress_module compress_230 (
                                            .x(u[0][230]),
                                            .d(10),
                                            .result(com_out[0][230])
                                        );
                                        
                                        compress_module compress_231 (
                                            .x(u[0][231]),
                                            .d(10),
                                            .result(com_out[0][231])
                                        );
                                        
                                        compress_module compress_232 (
                                            .x(u[0][232]),
                                            .d(10),
                                            .result(com_out[0][232])
                                        );
                                        
                                        compress_module compress_233 (
                                            .x(u[0][233]),
                                            .d(10),
                                            .result(com_out[0][233])
                                        );
                                        
                                        compress_module compress_234 (
                                            .x(u[0][234]),
                                            .d(10),
                                            .result(com_out[0][234])
                                        );
                                        
                                        compress_module compress_235 (
                                            .x(u[0][235]),
                                            .d(10),
                                            .result(com_out[0][235])
                                        );
                                        
                                        compress_module compress_236 (
                                            .x(u[0][236]),
                                            .d(10),
                                            .result(com_out[0][236])
                                        );
                                        
                                        compress_module compress_237 (
                                            .x(u[0][237]),
                                            .d(10),
                                            .result(com_out[0][237])
                                        );
                                        
                                        compress_module compress_238 (
                                            .x(u[0][238]),
                                            .d(10),
                                            .result(com_out[0][238])
                                        );
                                        
                                        compress_module compress_239 (
                                            .x(u[0][239]),
                                            .d(10),
                                            .result(com_out[0][239])
                                        );
                                        
                                        compress_module compress_240 (
                                            .x(u[0][240]),
                                            .d(10),
                                            .result(com_out[0][240])
                                        );
                                        
                                        compress_module compress_241 (
                                            .x(u[0][241]),
                                            .d(10),
                                            .result(com_out[0][241])
                                        );
                                        
                                        compress_module compress_242 (
                                            .x(u[0][242]),
                                            .d(10),
                                            .result(com_out[0][242])
                                        );
                                        
                                        compress_module compress_243 (
                                            .x(u[0][243]),
                                            .d(10),
                                            .result(com_out[0][243])
                                        );
                                        
                                        compress_module compress_244 (
                                            .x(u[0][244]),
                                            .d(10),
                                            .result(com_out[0][244])
                                        );
                                        
                                        compress_module compress_245 (
                                            .x(u[0][245]),
                                            .d(10),
                                            .result(com_out[0][245])
                                        );
                                        
                                        compress_module compress_246 (
                                            .x(u[0][246]),
                                            .d(10),
                                            .result(com_out[0][246])
                                        );
                                        
                                        compress_module compress_247 (
                                            .x(u[0][247]),
                                            .d(10),
                                            .result(com_out[0][247])
                                        );
                                        
                                        compress_module compress_248 (
                                            .x(u[0][248]),
                                            .d(10),
                                            .result(com_out[0][248])
                                        );
                                        
                                        compress_module compress_249 (
                                            .x(u[0][249]),
                                            .d(10),
                                            .result(com_out[0][249])
                                        );
                                        
                                        compress_module compress_250 (
                                            .x(u[0][250]),
                                            .d(10),
                                            .result(com_out[0][250])
                                        );
                                        
                                        compress_module compress_251 (
                                            .x(u[0][251]),
                                            .d(10),
                                            .result(com_out[0][251])
                                        );
                                        
                                        compress_module compress_252 (
                                            .x(u[0][252]),
                                            .d(10),
                                            .result(com_out[0][252])
                                        );
                                        
                                        compress_module compress_253 (
                                            .x(u[0][253]),
                                            .d(10),
                                            .result(com_out[0][253])
                                        );
                                        
                                        compress_module compress_254 (
                                            .x(u[0][254]),
                                            .d(10),
                                            .result(com_out[0][254])
                                        );
                                        
                                        compress_module compress_255 (
                                            .x(u[0][255]),
                                            .d(10),
                                            .result(com_out[0][255])
                                        );
                                        
                                        compress_module compress_256 (
                                            .x(u[1][0]),
                                            .d(10),
                                            .result(com_out[1][0])
                                        );
                                        
                                        compress_module compress_257 (
                                            .x(u[1][1]),
                                            .d(10),
                                            .result(com_out[1][1])
                                        );
                                        
                                        compress_module compress_258 (
                                            .x(u[1][2]),
                                            .d(10),
                                            .result(com_out[1][2])
                                        );
                                        
                                        compress_module compress_259 (
                                            .x(u[1][3]),
                                            .d(10),
                                            .result(com_out[1][3])
                                        );
                                        
                                        compress_module compress_260 (
                                            .x(u[1][4]),
                                            .d(10),
                                            .result(com_out[1][4])
                                        );
                                        
                                        compress_module compress_261 (
                                            .x(u[1][5]),
                                            .d(10),
                                            .result(com_out[1][5])
                                        );
                                        
                                        compress_module compress_262 (
                                            .x(u[1][6]),
                                            .d(10),
                                            .result(com_out[1][6])
                                        );
                                        
                                        compress_module compress_263 (
                                            .x(u[1][7]),
                                            .d(10),
                                            .result(com_out[1][7])
                                        );
                                        
                                        compress_module compress_264 (
                                            .x(u[1][8]),
                                            .d(10),
                                            .result(com_out[1][8])
                                        );
                                        
                                        compress_module compress_265 (
                                            .x(u[1][9]),
                                            .d(10),
                                            .result(com_out[1][9])
                                        );
                                        
                                        compress_module compress_266 (
                                            .x(u[1][10]),
                                            .d(10),
                                            .result(com_out[1][10])
                                        );
                                        
                                        compress_module compress_267 (
                                            .x(u[1][11]),
                                            .d(10),
                                            .result(com_out[1][11])
                                        );
                                        
                                        compress_module compress_268 (
                                            .x(u[1][12]),
                                            .d(10),
                                            .result(com_out[1][12])
                                        );
                                        
                                        compress_module compress_269 (
                                            .x(u[1][13]),
                                            .d(10),
                                            .result(com_out[1][13])
                                        );
                                        
                                        compress_module compress_270 (
                                            .x(u[1][14]),
                                            .d(10),
                                            .result(com_out[1][14])
                                        );
                                        
                                        compress_module compress_271 (
                                            .x(u[1][15]),
                                            .d(10),
                                            .result(com_out[1][15])
                                        );
                                        
                                        compress_module compress_272 (
                                            .x(u[1][16]),
                                            .d(10),
                                            .result(com_out[1][16])
                                        );
                                        
                                        compress_module compress_273 (
                                            .x(u[1][17]),
                                            .d(10),
                                            .result(com_out[1][17])
                                        );
                                        
                                        compress_module compress_274 (
                                            .x(u[1][18]),
                                            .d(10),
                                            .result(com_out[1][18])
                                        );
                                        
                                        compress_module compress_275 (
                                            .x(u[1][19]),
                                            .d(10),
                                            .result(com_out[1][19])
                                        );
                                        
                                        compress_module compress_276 (
                                            .x(u[1][20]),
                                            .d(10),
                                            .result(com_out[1][20])
                                        );
                                        
                                        compress_module compress_277 (
                                            .x(u[1][21]),
                                            .d(10),
                                            .result(com_out[1][21])
                                        );
                                        
                                        compress_module compress_278 (
                                            .x(u[1][22]),
                                            .d(10),
                                            .result(com_out[1][22])
                                        );
                                        
                                        compress_module compress_279 (
                                            .x(u[1][23]),
                                            .d(10),
                                            .result(com_out[1][23])
                                        );
                                        
                                        compress_module compress_280 (
                                            .x(u[1][24]),
                                            .d(10),
                                            .result(com_out[1][24])
                                        );
                                        
                                        compress_module compress_281 (
                                            .x(u[1][25]),
                                            .d(10),
                                            .result(com_out[1][25])
                                        );
                                        
                                        compress_module compress_282 (
                                            .x(u[1][26]),
                                            .d(10),
                                            .result(com_out[1][26])
                                        );
                                        
                                        compress_module compress_283 (
                                            .x(u[1][27]),
                                            .d(10),
                                            .result(com_out[1][27])
                                        );
                                        
                                        compress_module compress_284 (
                                            .x(u[1][28]),
                                            .d(10),
                                            .result(com_out[1][28])
                                        );
                                        
                                        compress_module compress_285 (
                                            .x(u[1][29]),
                                            .d(10),
                                            .result(com_out[1][29])
                                        );
                                        
                                        compress_module compress_286 (
                                            .x(u[1][30]),
                                            .d(10),
                                            .result(com_out[1][30])
                                        );
                                        
                                        compress_module compress_287 (
                                            .x(u[1][31]),
                                            .d(10),
                                            .result(com_out[1][31])
                                        );
                                        
                                        compress_module compress_288 (
                                            .x(u[1][32]),
                                            .d(10),
                                            .result(com_out[1][32])
                                        );
                                        
                                        compress_module compress_289 (
                                            .x(u[1][33]),
                                            .d(10),
                                            .result(com_out[1][33])
                                        );
                                        
                                        compress_module compress_290 (
                                            .x(u[1][34]),
                                            .d(10),
                                            .result(com_out[1][34])
                                        );
                                        
                                        compress_module compress_291 (
                                            .x(u[1][35]),
                                            .d(10),
                                            .result(com_out[1][35])
                                        );
                                        
                                        compress_module compress_292 (
                                            .x(u[1][36]),
                                            .d(10),
                                            .result(com_out[1][36])
                                        );
                                        
                                        compress_module compress_293 (
                                            .x(u[1][37]),
                                            .d(10),
                                            .result(com_out[1][37])
                                        );
                                        
                                        compress_module compress_294 (
                                            .x(u[1][38]),
                                            .d(10),
                                            .result(com_out[1][38])
                                        );
                                        
                                        compress_module compress_295 (
                                            .x(u[1][39]),
                                            .d(10),
                                            .result(com_out[1][39])
                                        );
                                        
                                        compress_module compress_296 (
                                            .x(u[1][40]),
                                            .d(10),
                                            .result(com_out[1][40])
                                        );
                                        
                                        compress_module compress_297 (
                                            .x(u[1][41]),
                                            .d(10),
                                            .result(com_out[1][41])
                                        );
                                        
                                        compress_module compress_298 (
                                            .x(u[1][42]),
                                            .d(10),
                                            .result(com_out[1][42])
                                        );
                                        
                                        compress_module compress_299 (
                                            .x(u[1][43]),
                                            .d(10),
                                            .result(com_out[1][43])
                                        );
                                        
                                        compress_module compress_300 (
                                            .x(u[1][44]),
                                            .d(10),
                                            .result(com_out[1][44])
                                        );
                                        
                                        compress_module compress_301 (
                                            .x(u[1][45]),
                                            .d(10),
                                            .result(com_out[1][45])
                                        );
                                        
                                        compress_module compress_302 (
                                            .x(u[1][46]),
                                            .d(10),
                                            .result(com_out[1][46])
                                        );
                                        
                                        compress_module compress_303 (
                                            .x(u[1][47]),
                                            .d(10),
                                            .result(com_out[1][47])
                                        );
                                        
                                        compress_module compress_304 (
                                            .x(u[1][48]),
                                            .d(10),
                                            .result(com_out[1][48])
                                        );
                                        
                                        compress_module compress_305 (
                                            .x(u[1][49]),
                                            .d(10),
                                            .result(com_out[1][49])
                                        );
                                        
                                        compress_module compress_306 (
                                            .x(u[1][50]),
                                            .d(10),
                                            .result(com_out[1][50])
                                        );
                                        
                                        compress_module compress_307 (
                                            .x(u[1][51]),
                                            .d(10),
                                            .result(com_out[1][51])
                                        );
                                        
                                        compress_module compress_308 (
                                            .x(u[1][52]),
                                            .d(10),
                                            .result(com_out[1][52])
                                        );
                                        
                                        compress_module compress_309 (
                                            .x(u[1][53]),
                                            .d(10),
                                            .result(com_out[1][53])
                                        );
                                        
                                        compress_module compress_310 (
                                            .x(u[1][54]),
                                            .d(10),
                                            .result(com_out[1][54])
                                        );
                                        
                                        compress_module compress_311 (
                                            .x(u[1][55]),
                                            .d(10),
                                            .result(com_out[1][55])
                                        );
                                        
                                        compress_module compress_312 (
                                            .x(u[1][56]),
                                            .d(10),
                                            .result(com_out[1][56])
                                        );
                                        
                                        compress_module compress_313 (
                                            .x(u[1][57]),
                                            .d(10),
                                            .result(com_out[1][57])
                                        );
                                        
                                        compress_module compress_314 (
                                            .x(u[1][58]),
                                            .d(10),
                                            .result(com_out[1][58])
                                        );
                                        
                                        compress_module compress_315 (
                                            .x(u[1][59]),
                                            .d(10),
                                            .result(com_out[1][59])
                                        );
                                        
                                        compress_module compress_316 (
                                            .x(u[1][60]),
                                            .d(10),
                                            .result(com_out[1][60])
                                        );
                                        
                                        compress_module compress_317 (
                                            .x(u[1][61]),
                                            .d(10),
                                            .result(com_out[1][61])
                                        );
                                        
                                        compress_module compress_318 (
                                            .x(u[1][62]),
                                            .d(10),
                                            .result(com_out[1][62])
                                        );
                                        
                                        compress_module compress_319 (
                                            .x(u[1][63]),
                                            .d(10),
                                            .result(com_out[1][63])
                                        );
                                        
                                        compress_module compress_320 (
                                            .x(u[1][64]),
                                            .d(10),
                                            .result(com_out[1][64])
                                        );
                                        
                                        compress_module compress_321 (
                                            .x(u[1][65]),
                                            .d(10),
                                            .result(com_out[1][65])
                                        );
                                        
                                        compress_module compress_322 (
                                            .x(u[1][66]),
                                            .d(10),
                                            .result(com_out[1][66])
                                        );
                                        
                                        compress_module compress_323 (
                                            .x(u[1][67]),
                                            .d(10),
                                            .result(com_out[1][67])
                                        );
                                        
                                        compress_module compress_324 (
                                            .x(u[1][68]),
                                            .d(10),
                                            .result(com_out[1][68])
                                        );
                                        
                                        compress_module compress_325 (
                                            .x(u[1][69]),
                                            .d(10),
                                            .result(com_out[1][69])
                                        );
                                        
                                        compress_module compress_326 (
                                            .x(u[1][70]),
                                            .d(10),
                                            .result(com_out[1][70])
                                        );
                                        
                                        compress_module compress_327 (
                                            .x(u[1][71]),
                                            .d(10),
                                            .result(com_out[1][71])
                                        );
                                        
                                        compress_module compress_328 (
                                            .x(u[1][72]),
                                            .d(10),
                                            .result(com_out[1][72])
                                        );
                                        
                                        compress_module compress_329 (
                                            .x(u[1][73]),
                                            .d(10),
                                            .result(com_out[1][73])
                                        );
                                        
                                        compress_module compress_330 (
                                            .x(u[1][74]),
                                            .d(10),
                                            .result(com_out[1][74])
                                        );
                                        
                                        compress_module compress_331 (
                                            .x(u[1][75]),
                                            .d(10),
                                            .result(com_out[1][75])
                                        );
                                        
                                        compress_module compress_332 (
                                            .x(u[1][76]),
                                            .d(10),
                                            .result(com_out[1][76])
                                        );
                                        
                                        compress_module compress_333 (
                                            .x(u[1][77]),
                                            .d(10),
                                            .result(com_out[1][77])
                                        );
                                        
                                        compress_module compress_334 (
                                            .x(u[1][78]),
                                            .d(10),
                                            .result(com_out[1][78])
                                        );
                                        
                                        compress_module compress_335 (
                                            .x(u[1][79]),
                                            .d(10),
                                            .result(com_out[1][79])
                                        );
                                        
                                        compress_module compress_336 (
                                            .x(u[1][80]),
                                            .d(10),
                                            .result(com_out[1][80])
                                        );
                                        
                                        compress_module compress_337 (
                                            .x(u[1][81]),
                                            .d(10),
                                            .result(com_out[1][81])
                                        );
                                        
                                        compress_module compress_338 (
                                            .x(u[1][82]),
                                            .d(10),
                                            .result(com_out[1][82])
                                        );
                                        
                                        compress_module compress_339 (
                                            .x(u[1][83]),
                                            .d(10),
                                            .result(com_out[1][83])
                                        );
                                        
                                        compress_module compress_340 (
                                            .x(u[1][84]),
                                            .d(10),
                                            .result(com_out[1][84])
                                        );
                                        
                                        compress_module compress_341 (
                                            .x(u[1][85]),
                                            .d(10),
                                            .result(com_out[1][85])
                                        );
                                        
                                        compress_module compress_342 (
                                            .x(u[1][86]),
                                            .d(10),
                                            .result(com_out[1][86])
                                        );
                                        
                                        compress_module compress_343 (
                                            .x(u[1][87]),
                                            .d(10),
                                            .result(com_out[1][87])
                                        );
                                        
                                        compress_module compress_344 (
                                            .x(u[1][88]),
                                            .d(10),
                                            .result(com_out[1][88])
                                        );
                                        
                                        compress_module compress_345 (
                                            .x(u[1][89]),
                                            .d(10),
                                            .result(com_out[1][89])
                                        );
                                        
                                        compress_module compress_346 (
                                            .x(u[1][90]),
                                            .d(10),
                                            .result(com_out[1][90])
                                        );
                                        
                                        compress_module compress_347 (
                                            .x(u[1][91]),
                                            .d(10),
                                            .result(com_out[1][91])
                                        );
                                        
                                        compress_module compress_348 (
                                            .x(u[1][92]),
                                            .d(10),
                                            .result(com_out[1][92])
                                        );
                                        
                                        compress_module compress_349 (
                                            .x(u[1][93]),
                                            .d(10),
                                            .result(com_out[1][93])
                                        );
                                        
                                        compress_module compress_350 (
                                            .x(u[1][94]),
                                            .d(10),
                                            .result(com_out[1][94])
                                        );
                                        
                                        compress_module compress_351 (
                                            .x(u[1][95]),
                                            .d(10),
                                            .result(com_out[1][95])
                                        );
                                        
                                        compress_module compress_352 (
                                            .x(u[1][96]),
                                            .d(10),
                                            .result(com_out[1][96])
                                        );
                                        
                                        compress_module compress_353 (
                                            .x(u[1][97]),
                                            .d(10),
                                            .result(com_out[1][97])
                                        );
                                        
                                        compress_module compress_354 (
                                            .x(u[1][98]),
                                            .d(10),
                                            .result(com_out[1][98])
                                        );
                                        
                                        compress_module compress_355 (
                                            .x(u[1][99]),
                                            .d(10),
                                            .result(com_out[1][99])
                                        );
                                        
                                        compress_module compress_356 (
                                            .x(u[1][100]),
                                            .d(10),
                                            .result(com_out[1][100])
                                        );
                                        
                                        compress_module compress_357 (
                                            .x(u[1][101]),
                                            .d(10),
                                            .result(com_out[1][101])
                                        );
                                        
                                        compress_module compress_358 (
                                            .x(u[1][102]),
                                            .d(10),
                                            .result(com_out[1][102])
                                        );
                                        
                                        compress_module compress_359 (
                                            .x(u[1][103]),
                                            .d(10),
                                            .result(com_out[1][103])
                                        );
                                        
                                        compress_module compress_360 (
                                            .x(u[1][104]),
                                            .d(10),
                                            .result(com_out[1][104])
                                        );
                                        
                                        compress_module compress_361 (
                                            .x(u[1][105]),
                                            .d(10),
                                            .result(com_out[1][105])
                                        );
                                        
                                        compress_module compress_362 (
                                            .x(u[1][106]),
                                            .d(10),
                                            .result(com_out[1][106])
                                        );
                                        
                                        compress_module compress_363 (
                                            .x(u[1][107]),
                                            .d(10),
                                            .result(com_out[1][107])
                                        );
                                        
                                        compress_module compress_364 (
                                            .x(u[1][108]),
                                            .d(10),
                                            .result(com_out[1][108])
                                        );
                                        
                                        compress_module compress_365 (
                                            .x(u[1][109]),
                                            .d(10),
                                            .result(com_out[1][109])
                                        );
                                        
                                        compress_module compress_366 (
                                            .x(u[1][110]),
                                            .d(10),
                                            .result(com_out[1][110])
                                        );
                                        
                                        compress_module compress_367 (
                                            .x(u[1][111]),
                                            .d(10),
                                            .result(com_out[1][111])
                                        );
                                        
                                        compress_module compress_368 (
                                            .x(u[1][112]),
                                            .d(10),
                                            .result(com_out[1][112])
                                        );
                                        
                                        compress_module compress_369 (
                                            .x(u[1][113]),
                                            .d(10),
                                            .result(com_out[1][113])
                                        );
                                        
                                        compress_module compress_370 (
                                            .x(u[1][114]),
                                            .d(10),
                                            .result(com_out[1][114])
                                        );
                                        
                                        compress_module compress_371 (
                                            .x(u[1][115]),
                                            .d(10),
                                            .result(com_out[1][115])
                                        );
                                        
                                        compress_module compress_372 (
                                            .x(u[1][116]),
                                            .d(10),
                                            .result(com_out[1][116])
                                        );
                                        
                                        compress_module compress_373 (
                                            .x(u[1][117]),
                                            .d(10),
                                            .result(com_out[1][117])
                                        );
                                        
                                        compress_module compress_374 (
                                            .x(u[1][118]),
                                            .d(10),
                                            .result(com_out[1][118])
                                        );
                                        
                                        compress_module compress_375 (
                                            .x(u[1][119]),
                                            .d(10),
                                            .result(com_out[1][119])
                                        );
                                        
                                        compress_module compress_376 (
                                            .x(u[1][120]),
                                            .d(10),
                                            .result(com_out[1][120])
                                        );
                                        
                                        compress_module compress_377 (
                                            .x(u[1][121]),
                                            .d(10),
                                            .result(com_out[1][121])
                                        );
                                        
                                        compress_module compress_378 (
                                            .x(u[1][122]),
                                            .d(10),
                                            .result(com_out[1][122])
                                        );
                                        
                                        compress_module compress_379 (
                                            .x(u[1][123]),
                                            .d(10),
                                            .result(com_out[1][123])
                                        );
                                        
                                        compress_module compress_380 (
                                            .x(u[1][124]),
                                            .d(10),
                                            .result(com_out[1][124])
                                        );
                                        
                                        compress_module compress_381 (
                                            .x(u[1][125]),
                                            .d(10),
                                            .result(com_out[1][125])
                                        );
                                        
                                        compress_module compress_382 (
                                            .x(u[1][126]),
                                            .d(10),
                                            .result(com_out[1][126])
                                        );
                                        
                                        compress_module compress_383 (
                                            .x(u[1][127]),
                                            .d(10),
                                            .result(com_out[1][127])
                                        );
                                        
                                        compress_module compress_384 (
                                            .x(u[1][128]),
                                            .d(10),
                                            .result(com_out[1][128])
                                        );
                                        
                                        compress_module compress_385 (
                                            .x(u[1][129]),
                                            .d(10),
                                            .result(com_out[1][129])
                                        );
                                        
                                        compress_module compress_386 (
                                            .x(u[1][130]),
                                            .d(10),
                                            .result(com_out[1][130])
                                        );
                                        
                                        compress_module compress_387 (
                                            .x(u[1][131]),
                                            .d(10),
                                            .result(com_out[1][131])
                                        );
                                        
                                        compress_module compress_388 (
                                            .x(u[1][132]),
                                            .d(10),
                                            .result(com_out[1][132])
                                        );
                                        
                                        compress_module compress_389 (
                                            .x(u[1][133]),
                                            .d(10),
                                            .result(com_out[1][133])
                                        );
                                        
                                        compress_module compress_390 (
                                            .x(u[1][134]),
                                            .d(10),
                                            .result(com_out[1][134])
                                        );
                                        
                                        compress_module compress_391 (
                                            .x(u[1][135]),
                                            .d(10),
                                            .result(com_out[1][135])
                                        );
                                        
                                        compress_module compress_392 (
                                            .x(u[1][136]),
                                            .d(10),
                                            .result(com_out[1][136])
                                        );
                                        
                                        compress_module compress_393 (
                                            .x(u[1][137]),
                                            .d(10),
                                            .result(com_out[1][137])
                                        );
                                        
                                        compress_module compress_394 (
                                            .x(u[1][138]),
                                            .d(10),
                                            .result(com_out[1][138])
                                        );
                                        
                                        compress_module compress_395 (
                                            .x(u[1][139]),
                                            .d(10),
                                            .result(com_out[1][139])
                                        );
                                        
                                        compress_module compress_396 (
                                            .x(u[1][140]),
                                            .d(10),
                                            .result(com_out[1][140])
                                        );
                                        
                                        compress_module compress_397 (
                                            .x(u[1][141]),
                                            .d(10),
                                            .result(com_out[1][141])
                                        );
                                        
                                        compress_module compress_398 (
                                            .x(u[1][142]),
                                            .d(10),
                                            .result(com_out[1][142])
                                        );
                                        
                                        compress_module compress_399 (
                                            .x(u[1][143]),
                                            .d(10),
                                            .result(com_out[1][143])
                                        );
                                        
                                        compress_module compress_400 (
                                            .x(u[1][144]),
                                            .d(10),
                                            .result(com_out[1][144])
                                        );
                                        
                                        compress_module compress_401 (
                                            .x(u[1][145]),
                                            .d(10),
                                            .result(com_out[1][145])
                                        );
                                        
                                        compress_module compress_402 (
                                            .x(u[1][146]),
                                            .d(10),
                                            .result(com_out[1][146])
                                        );
                                        
                                        compress_module compress_403 (
                                            .x(u[1][147]),
                                            .d(10),
                                            .result(com_out[1][147])
                                        );
                                        
                                        compress_module compress_404 (
                                            .x(u[1][148]),
                                            .d(10),
                                            .result(com_out[1][148])
                                        );
                                        
                                        compress_module compress_405 (
                                            .x(u[1][149]),
                                            .d(10),
                                            .result(com_out[1][149])
                                        );
                                        
                                        compress_module compress_406 (
                                            .x(u[1][150]),
                                            .d(10),
                                            .result(com_out[1][150])
                                        );
                                        
                                        compress_module compress_407 (
                                            .x(u[1][151]),
                                            .d(10),
                                            .result(com_out[1][151])
                                        );
                                        
                                        compress_module compress_408 (
                                            .x(u[1][152]),
                                            .d(10),
                                            .result(com_out[1][152])
                                        );
                                        
                                        compress_module compress_409 (
                                            .x(u[1][153]),
                                            .d(10),
                                            .result(com_out[1][153])
                                        );
                                        
                                        compress_module compress_410 (
                                            .x(u[1][154]),
                                            .d(10),
                                            .result(com_out[1][154])
                                        );
                                        
                                        compress_module compress_411 (
                                            .x(u[1][155]),
                                            .d(10),
                                            .result(com_out[1][155])
                                        );
                                        
                                        compress_module compress_412 (
                                            .x(u[1][156]),
                                            .d(10),
                                            .result(com_out[1][156])
                                        );
                                        
                                        compress_module compress_413 (
                                            .x(u[1][157]),
                                            .d(10),
                                            .result(com_out[1][157])
                                        );
                                        
                                        compress_module compress_414 (
                                            .x(u[1][158]),
                                            .d(10),
                                            .result(com_out[1][158])
                                        );
                                        
                                        compress_module compress_415 (
                                            .x(u[1][159]),
                                            .d(10),
                                            .result(com_out[1][159])
                                        );
                                        
                                        compress_module compress_416 (
                                            .x(u[1][160]),
                                            .d(10),
                                            .result(com_out[1][160])
                                        );
                                        
                                        compress_module compress_417 (
                                            .x(u[1][161]),
                                            .d(10),
                                            .result(com_out[1][161])
                                        );
                                        
                                        compress_module compress_418 (
                                            .x(u[1][162]),
                                            .d(10),
                                            .result(com_out[1][162])
                                        );
                                        
                                        compress_module compress_419 (
                                            .x(u[1][163]),
                                            .d(10),
                                            .result(com_out[1][163])
                                        );
                                        
                                        compress_module compress_420 (
                                            .x(u[1][164]),
                                            .d(10),
                                            .result(com_out[1][164])
                                        );
                                        
                                        compress_module compress_421 (
                                            .x(u[1][165]),
                                            .d(10),
                                            .result(com_out[1][165])
                                        );
                                        
                                        compress_module compress_422 (
                                            .x(u[1][166]),
                                            .d(10),
                                            .result(com_out[1][166])
                                        );
                                        
                                        compress_module compress_423 (
                                            .x(u[1][167]),
                                            .d(10),
                                            .result(com_out[1][167])
                                        );
                                        
                                        compress_module compress_424 (
                                            .x(u[1][168]),
                                            .d(10),
                                            .result(com_out[1][168])
                                        );
                                        
                                        compress_module compress_425 (
                                            .x(u[1][169]),
                                            .d(10),
                                            .result(com_out[1][169])
                                        );
                                        
                                        compress_module compress_426 (
                                            .x(u[1][170]),
                                            .d(10),
                                            .result(com_out[1][170])
                                        );
                                        
                                        compress_module compress_427 (
                                            .x(u[1][171]),
                                            .d(10),
                                            .result(com_out[1][171])
                                        );
                                        
                                        compress_module compress_428 (
                                            .x(u[1][172]),
                                            .d(10),
                                            .result(com_out[1][172])
                                        );
                                        
                                        compress_module compress_429 (
                                            .x(u[1][173]),
                                            .d(10),
                                            .result(com_out[1][173])
                                        );
                                        
                                        compress_module compress_430 (
                                            .x(u[1][174]),
                                            .d(10),
                                            .result(com_out[1][174])
                                        );
                                        
                                        compress_module compress_431 (
                                            .x(u[1][175]),
                                            .d(10),
                                            .result(com_out[1][175])
                                        );
                                        
                                        compress_module compress_432 (
                                            .x(u[1][176]),
                                            .d(10),
                                            .result(com_out[1][176])
                                        );
                                        
                                        compress_module compress_433 (
                                            .x(u[1][177]),
                                            .d(10),
                                            .result(com_out[1][177])
                                        );
                                        
                                        compress_module compress_434 (
                                            .x(u[1][178]),
                                            .d(10),
                                            .result(com_out[1][178])
                                        );
                                        
                                        compress_module compress_435 (
                                            .x(u[1][179]),
                                            .d(10),
                                            .result(com_out[1][179])
                                        );
                                        
                                        compress_module compress_436 (
                                            .x(u[1][180]),
                                            .d(10),
                                            .result(com_out[1][180])
                                        );
                                        
                                        compress_module compress_437 (
                                            .x(u[1][181]),
                                            .d(10),
                                            .result(com_out[1][181])
                                        );
                                        
                                        compress_module compress_438 (
                                            .x(u[1][182]),
                                            .d(10),
                                            .result(com_out[1][182])
                                        );
                                        
                                        compress_module compress_439 (
                                            .x(u[1][183]),
                                            .d(10),
                                            .result(com_out[1][183])
                                        );
                                        
                                        compress_module compress_440 (
                                            .x(u[1][184]),
                                            .d(10),
                                            .result(com_out[1][184])
                                        );
                                        
                                        compress_module compress_441 (
                                            .x(u[1][185]),
                                            .d(10),
                                            .result(com_out[1][185])
                                        );
                                        
                                        compress_module compress_442 (
                                            .x(u[1][186]),
                                            .d(10),
                                            .result(com_out[1][186])
                                        );
                                        
                                        compress_module compress_443 (
                                            .x(u[1][187]),
                                            .d(10),
                                            .result(com_out[1][187])
                                        );
                                        
                                        compress_module compress_444 (
                                            .x(u[1][188]),
                                            .d(10),
                                            .result(com_out[1][188])
                                        );
                                        
                                        compress_module compress_445 (
                                            .x(u[1][189]),
                                            .d(10),
                                            .result(com_out[1][189])
                                        );
                                        
                                        compress_module compress_446 (
                                            .x(u[1][190]),
                                            .d(10),
                                            .result(com_out[1][190])
                                        );
                                        
                                        compress_module compress_447 (
                                            .x(u[1][191]),
                                            .d(10),
                                            .result(com_out[1][191])
                                        );
                                        
                                        compress_module compress_448 (
                                            .x(u[1][192]),
                                            .d(10),
                                            .result(com_out[1][192])
                                        );
                                        
                                        compress_module compress_449 (
                                            .x(u[1][193]),
                                            .d(10),
                                            .result(com_out[1][193])
                                        );
                                        
                                        compress_module compress_450 (
                                            .x(u[1][194]),
                                            .d(10),
                                            .result(com_out[1][194])
                                        );
                                        
                                        compress_module compress_451 (
                                            .x(u[1][195]),
                                            .d(10),
                                            .result(com_out[1][195])
                                        );
                                        
                                        compress_module compress_452 (
                                            .x(u[1][196]),
                                            .d(10),
                                            .result(com_out[1][196])
                                        );
                                        
                                        compress_module compress_453 (
                                            .x(u[1][197]),
                                            .d(10),
                                            .result(com_out[1][197])
                                        );
                                        
                                        compress_module compress_454 (
                                            .x(u[1][198]),
                                            .d(10),
                                            .result(com_out[1][198])
                                        );
                                        
                                        compress_module compress_455 (
                                            .x(u[1][199]),
                                            .d(10),
                                            .result(com_out[1][199])
                                        );
                                        
                                        compress_module compress_456 (
                                            .x(u[1][200]),
                                            .d(10),
                                            .result(com_out[1][200])
                                        );
                                        
                                        compress_module compress_457 (
                                            .x(u[1][201]),
                                            .d(10),
                                            .result(com_out[1][201])
                                        );
                                        
                                        compress_module compress_458 (
                                            .x(u[1][202]),
                                            .d(10),
                                            .result(com_out[1][202])
                                        );
                                        
                                        compress_module compress_459 (
                                            .x(u[1][203]),
                                            .d(10),
                                            .result(com_out[1][203])
                                        );
                                        
                                        compress_module compress_460 (
                                            .x(u[1][204]),
                                            .d(10),
                                            .result(com_out[1][204])
                                        );
                                        
                                        compress_module compress_461 (
                                            .x(u[1][205]),
                                            .d(10),
                                            .result(com_out[1][205])
                                        );
                                        
                                        compress_module compress_462 (
                                            .x(u[1][206]),
                                            .d(10),
                                            .result(com_out[1][206])
                                        );
                                        
                                        compress_module compress_463 (
                                            .x(u[1][207]),
                                            .d(10),
                                            .result(com_out[1][207])
                                        );
                                        
                                        compress_module compress_464 (
                                            .x(u[1][208]),
                                            .d(10),
                                            .result(com_out[1][208])
                                        );
                                        
                                        compress_module compress_465 (
                                            .x(u[1][209]),
                                            .d(10),
                                            .result(com_out[1][209])
                                        );
                                        
                                        compress_module compress_466 (
                                            .x(u[1][210]),
                                            .d(10),
                                            .result(com_out[1][210])
                                        );
                                        
                                        compress_module compress_467 (
                                            .x(u[1][211]),
                                            .d(10),
                                            .result(com_out[1][211])
                                        );
                                        
                                        compress_module compress_468 (
                                            .x(u[1][212]),
                                            .d(10),
                                            .result(com_out[1][212])
                                        );
                                        
                                        compress_module compress_469 (
                                            .x(u[1][213]),
                                            .d(10),
                                            .result(com_out[1][213])
                                        );
                                        
                                        compress_module compress_470 (
                                            .x(u[1][214]),
                                            .d(10),
                                            .result(com_out[1][214])
                                        );
                                        
                                        compress_module compress_471 (
                                            .x(u[1][215]),
                                            .d(10),
                                            .result(com_out[1][215])
                                        );
                                        
                                        compress_module compress_472 (
                                            .x(u[1][216]),
                                            .d(10),
                                            .result(com_out[1][216])
                                        );
                                        
                                        compress_module compress_473 (
                                            .x(u[1][217]),
                                            .d(10),
                                            .result(com_out[1][217])
                                        );
                                        
                                        compress_module compress_474 (
                                            .x(u[1][218]),
                                            .d(10),
                                            .result(com_out[1][218])
                                        );
                                        
                                        compress_module compress_475 (
                                            .x(u[1][219]),
                                            .d(10),
                                            .result(com_out[1][219])
                                        );
                                        
                                        compress_module compress_476 (
                                            .x(u[1][220]),
                                            .d(10),
                                            .result(com_out[1][220])
                                        );
                                        
                                        compress_module compress_477 (
                                            .x(u[1][221]),
                                            .d(10),
                                            .result(com_out[1][221])
                                        );
                                        
                                        compress_module compress_478 (
                                            .x(u[1][222]),
                                            .d(10),
                                            .result(com_out[1][222])
                                        );
                                        
                                        compress_module compress_479 (
                                            .x(u[1][223]),
                                            .d(10),
                                            .result(com_out[1][223])
                                        );
                                        
                                        compress_module compress_480 (
                                            .x(u[1][224]),
                                            .d(10),
                                            .result(com_out[1][224])
                                        );
                                        
                                        compress_module compress_481 (
                                            .x(u[1][225]),
                                            .d(10),
                                            .result(com_out[1][225])
                                        );
                                        
                                        compress_module compress_482 (
                                            .x(u[1][226]),
                                            .d(10),
                                            .result(com_out[1][226])
                                        );
                                        
                                        compress_module compress_483 (
                                            .x(u[1][227]),
                                            .d(10),
                                            .result(com_out[1][227])
                                        );
                                        
                                        compress_module compress_484 (
                                            .x(u[1][228]),
                                            .d(10),
                                            .result(com_out[1][228])
                                        );
                                        
                                        compress_module compress_485 (
                                            .x(u[1][229]),
                                            .d(10),
                                            .result(com_out[1][229])
                                        );
                                        
                                        compress_module compress_486 (
                                            .x(u[1][230]),
                                            .d(10),
                                            .result(com_out[1][230])
                                        );
                                        
                                        compress_module compress_487 (
                                            .x(u[1][231]),
                                            .d(10),
                                            .result(com_out[1][231])
                                        );
                                        
                                        compress_module compress_488 (
                                            .x(u[1][232]),
                                            .d(10),
                                            .result(com_out[1][232])
                                        );
                                        
                                        compress_module compress_489 (
                                            .x(u[1][233]),
                                            .d(10),
                                            .result(com_out[1][233])
                                        );
                                        
                                        compress_module compress_490 (
                                            .x(u[1][234]),
                                            .d(10),
                                            .result(com_out[1][234])
                                        );
                                        
                                        compress_module compress_491 (
                                            .x(u[1][235]),
                                            .d(10),
                                            .result(com_out[1][235])
                                        );
                                        
                                        compress_module compress_492 (
                                            .x(u[1][236]),
                                            .d(10),
                                            .result(com_out[1][236])
                                        );
                                        
                                        compress_module compress_493 (
                                            .x(u[1][237]),
                                            .d(10),
                                            .result(com_out[1][237])
                                        );
                                        
                                        compress_module compress_494 (
                                            .x(u[1][238]),
                                            .d(10),
                                            .result(com_out[1][238])
                                        );
                                        
                                        compress_module compress_495 (
                                            .x(u[1][239]),
                                            .d(10),
                                            .result(com_out[1][239])
                                        );
                                        
                                        compress_module compress_496 (
                                            .x(u[1][240]),
                                            .d(10),
                                            .result(com_out[1][240])
                                        );
                                        
                                        compress_module compress_497 (
                                            .x(u[1][241]),
                                            .d(10),
                                            .result(com_out[1][241])
                                        );
                                        
                                        compress_module compress_498 (
                                            .x(u[1][242]),
                                            .d(10),
                                            .result(com_out[1][242])
                                        );
                                        
                                        compress_module compress_499 (
                                            .x(u[1][243]),
                                            .d(10),
                                            .result(com_out[1][243])
                                        );
                                        
                                        compress_module compress_500 (
                                            .x(u[1][244]),
                                            .d(10),
                                            .result(com_out[1][244])
                                        );
                                        
                                        compress_module compress_501 (
                                            .x(u[1][245]),
                                            .d(10),
                                            .result(com_out[1][245])
                                        );
                                        
                                        compress_module compress_502 (
                                            .x(u[1][246]),
                                            .d(10),
                                            .result(com_out[1][246])
                                        );
                                        
                                        compress_module compress_503 (
                                            .x(u[1][247]),
                                            .d(10),
                                            .result(com_out[1][247])
                                        );
                                        
                                        compress_module compress_504 (
                                            .x(u[1][248]),
                                            .d(10),
                                            .result(com_out[1][248])
                                        );
                                        
                                        compress_module compress_505 (
                                            .x(u[1][249]),
                                            .d(10),
                                            .result(com_out[1][249])
                                        );
                                        
                                        compress_module compress_506 (
                                            .x(u[1][250]),
                                            .d(10),
                                            .result(com_out[1][250])
                                        );
                                        
                                        compress_module compress_507 (
                                            .x(u[1][251]),
                                            .d(10),
                                            .result(com_out[1][251])
                                        );
                                        
                                        compress_module compress_508 (
                                            .x(u[1][252]),
                                            .d(10),
                                            .result(com_out[1][252])
                                        );
                                        
                                        compress_module compress_509 (
                                            .x(u[1][253]),
                                            .d(10),
                                            .result(com_out[1][253])
                                        );
                                        
                                        compress_module compress_510 (
                                            .x(u[1][254]),
                                            .d(10),
                                            .result(com_out[1][254])
                                        );
                                        
                                        compress_module compress_511 (
                                            .x(u[1][255]),
                                            .d(10),
                                            .result(com_out[1][255])
                                        );
                                        
                                        compress_module compress_512 (
                                            .x(u[2][0]),
                                            .d(10),
                                            .result(com_out[2][0])
                                        );
                                        
                                        compress_module compress_513 (
                                            .x(u[2][1]),
                                            .d(10),
                                            .result(com_out[2][1])
                                        );
                                        
                                        compress_module compress_514 (
                                            .x(u[2][2]),
                                            .d(10),
                                            .result(com_out[2][2])
                                        );
                                        
                                        compress_module compress_515 (
                                            .x(u[2][3]),
                                            .d(10),
                                            .result(com_out[2][3])
                                        );
                                        
                                        compress_module compress_516 (
                                            .x(u[2][4]),
                                            .d(10),
                                            .result(com_out[2][4])
                                        );
                                        
                                        compress_module compress_517 (
                                            .x(u[2][5]),
                                            .d(10),
                                            .result(com_out[2][5])
                                        );
                                        
                                        compress_module compress_518 (
                                            .x(u[2][6]),
                                            .d(10),
                                            .result(com_out[2][6])
                                        );
                                        
                                        compress_module compress_519 (
                                            .x(u[2][7]),
                                            .d(10),
                                            .result(com_out[2][7])
                                        );
                                        
                                        compress_module compress_520 (
                                            .x(u[2][8]),
                                            .d(10),
                                            .result(com_out[2][8])
                                        );
                                        
                                        compress_module compress_521 (
                                            .x(u[2][9]),
                                            .d(10),
                                            .result(com_out[2][9])
                                        );
                                        
                                        compress_module compress_522 (
                                            .x(u[2][10]),
                                            .d(10),
                                            .result(com_out[2][10])
                                        );
                                        
                                        compress_module compress_523 (
                                            .x(u[2][11]),
                                            .d(10),
                                            .result(com_out[2][11])
                                        );
                                        
                                        compress_module compress_524 (
                                            .x(u[2][12]),
                                            .d(10),
                                            .result(com_out[2][12])
                                        );
                                        
                                        compress_module compress_525 (
                                            .x(u[2][13]),
                                            .d(10),
                                            .result(com_out[2][13])
                                        );
                                        
                                        compress_module compress_526 (
                                            .x(u[2][14]),
                                            .d(10),
                                            .result(com_out[2][14])
                                        );
                                        
                                        compress_module compress_527 (
                                            .x(u[2][15]),
                                            .d(10),
                                            .result(com_out[2][15])
                                        );
                                        
                                        compress_module compress_528 (
                                            .x(u[2][16]),
                                            .d(10),
                                            .result(com_out[2][16])
                                        );
                                        
                                        compress_module compress_529 (
                                            .x(u[2][17]),
                                            .d(10),
                                            .result(com_out[2][17])
                                        );
                                        
                                        compress_module compress_530 (
                                            .x(u[2][18]),
                                            .d(10),
                                            .result(com_out[2][18])
                                        );
                                        
                                        compress_module compress_531 (
                                            .x(u[2][19]),
                                            .d(10),
                                            .result(com_out[2][19])
                                        );
                                        
                                        compress_module compress_532 (
                                            .x(u[2][20]),
                                            .d(10),
                                            .result(com_out[2][20])
                                        );
                                        
                                        compress_module compress_533 (
                                            .x(u[2][21]),
                                            .d(10),
                                            .result(com_out[2][21])
                                        );
                                        
                                        compress_module compress_534 (
                                            .x(u[2][22]),
                                            .d(10),
                                            .result(com_out[2][22])
                                        );
                                        
                                        compress_module compress_535 (
                                            .x(u[2][23]),
                                            .d(10),
                                            .result(com_out[2][23])
                                        );
                                        
                                        compress_module compress_536 (
                                            .x(u[2][24]),
                                            .d(10),
                                            .result(com_out[2][24])
                                        );
                                        
                                        compress_module compress_537 (
                                            .x(u[2][25]),
                                            .d(10),
                                            .result(com_out[2][25])
                                        );
                                        
                                        compress_module compress_538 (
                                            .x(u[2][26]),
                                            .d(10),
                                            .result(com_out[2][26])
                                        );
                                        
                                        compress_module compress_539 (
                                            .x(u[2][27]),
                                            .d(10),
                                            .result(com_out[2][27])
                                        );
                                        
                                        compress_module compress_540 (
                                            .x(u[2][28]),
                                            .d(10),
                                            .result(com_out[2][28])
                                        );
                                        
                                        compress_module compress_541 (
                                            .x(u[2][29]),
                                            .d(10),
                                            .result(com_out[2][29])
                                        );
                                        
                                        compress_module compress_542 (
                                            .x(u[2][30]),
                                            .d(10),
                                            .result(com_out[2][30])
                                        );
                                        
                                        compress_module compress_543 (
                                            .x(u[2][31]),
                                            .d(10),
                                            .result(com_out[2][31])
                                        );
                                        
                                        compress_module compress_544 (
                                            .x(u[2][32]),
                                            .d(10),
                                            .result(com_out[2][32])
                                        );
                                        
                                        compress_module compress_545 (
                                            .x(u[2][33]),
                                            .d(10),
                                            .result(com_out[2][33])
                                        );
                                        
                                        compress_module compress_546 (
                                            .x(u[2][34]),
                                            .d(10),
                                            .result(com_out[2][34])
                                        );
                                        
                                        compress_module compress_547 (
                                            .x(u[2][35]),
                                            .d(10),
                                            .result(com_out[2][35])
                                        );
                                        
                                        compress_module compress_548 (
                                            .x(u[2][36]),
                                            .d(10),
                                            .result(com_out[2][36])
                                        );
                                        
                                        compress_module compress_549 (
                                            .x(u[2][37]),
                                            .d(10),
                                            .result(com_out[2][37])
                                        );
                                        
                                        compress_module compress_550 (
                                            .x(u[2][38]),
                                            .d(10),
                                            .result(com_out[2][38])
                                        );
                                        
                                        compress_module compress_551 (
                                            .x(u[2][39]),
                                            .d(10),
                                            .result(com_out[2][39])
                                        );
                                        
                                        compress_module compress_552 (
                                            .x(u[2][40]),
                                            .d(10),
                                            .result(com_out[2][40])
                                        );
                                        
                                        compress_module compress_553 (
                                            .x(u[2][41]),
                                            .d(10),
                                            .result(com_out[2][41])
                                        );
                                        
                                        compress_module compress_554 (
                                            .x(u[2][42]),
                                            .d(10),
                                            .result(com_out[2][42])
                                        );
                                        
                                        compress_module compress_555 (
                                            .x(u[2][43]),
                                            .d(10),
                                            .result(com_out[2][43])
                                        );
                                        
                                        compress_module compress_556 (
                                            .x(u[2][44]),
                                            .d(10),
                                            .result(com_out[2][44])
                                        );
                                        
                                        compress_module compress_557 (
                                            .x(u[2][45]),
                                            .d(10),
                                            .result(com_out[2][45])
                                        );
                                        
                                        compress_module compress_558 (
                                            .x(u[2][46]),
                                            .d(10),
                                            .result(com_out[2][46])
                                        );
                                        
                                        compress_module compress_559 (
                                            .x(u[2][47]),
                                            .d(10),
                                            .result(com_out[2][47])
                                        );
                                        
                                        compress_module compress_560 (
                                            .x(u[2][48]),
                                            .d(10),
                                            .result(com_out[2][48])
                                        );
                                        
                                        compress_module compress_561 (
                                            .x(u[2][49]),
                                            .d(10),
                                            .result(com_out[2][49])
                                        );
                                        
                                        compress_module compress_562 (
                                            .x(u[2][50]),
                                            .d(10),
                                            .result(com_out[2][50])
                                        );
                                        
                                        compress_module compress_563 (
                                            .x(u[2][51]),
                                            .d(10),
                                            .result(com_out[2][51])
                                        );
                                        
                                        compress_module compress_564 (
                                            .x(u[2][52]),
                                            .d(10),
                                            .result(com_out[2][52])
                                        );
                                        
                                        compress_module compress_565 (
                                            .x(u[2][53]),
                                            .d(10),
                                            .result(com_out[2][53])
                                        );
                                        
                                        compress_module compress_566 (
                                            .x(u[2][54]),
                                            .d(10),
                                            .result(com_out[2][54])
                                        );
                                        
                                        compress_module compress_567 (
                                            .x(u[2][55]),
                                            .d(10),
                                            .result(com_out[2][55])
                                        );
                                        
                                        compress_module compress_568 (
                                            .x(u[2][56]),
                                            .d(10),
                                            .result(com_out[2][56])
                                        );
                                        
                                        compress_module compress_569 (
                                            .x(u[2][57]),
                                            .d(10),
                                            .result(com_out[2][57])
                                        );
                                        
                                        compress_module compress_570 (
                                            .x(u[2][58]),
                                            .d(10),
                                            .result(com_out[2][58])
                                        );
                                        
                                        compress_module compress_571 (
                                            .x(u[2][59]),
                                            .d(10),
                                            .result(com_out[2][59])
                                        );
                                        
                                        compress_module compress_572 (
                                            .x(u[2][60]),
                                            .d(10),
                                            .result(com_out[2][60])
                                        );
                                        
                                        compress_module compress_573 (
                                            .x(u[2][61]),
                                            .d(10),
                                            .result(com_out[2][61])
                                        );
                                        
                                        compress_module compress_574 (
                                            .x(u[2][62]),
                                            .d(10),
                                            .result(com_out[2][62])
                                        );
                                        
                                        compress_module compress_575 (
                                            .x(u[2][63]),
                                            .d(10),
                                            .result(com_out[2][63])
                                        );
                                        
                                        compress_module compress_576 (
                                            .x(u[2][64]),
                                            .d(10),
                                            .result(com_out[2][64])
                                        );
                                        
                                        compress_module compress_577 (
                                            .x(u[2][65]),
                                            .d(10),
                                            .result(com_out[2][65])
                                        );
                                        
                                        compress_module compress_578 (
                                            .x(u[2][66]),
                                            .d(10),
                                            .result(com_out[2][66])
                                        );
                                        
                                        compress_module compress_579 (
                                            .x(u[2][67]),
                                            .d(10),
                                            .result(com_out[2][67])
                                        );
                                        
                                        compress_module compress_580 (
                                            .x(u[2][68]),
                                            .d(10),
                                            .result(com_out[2][68])
                                        );
                                        
                                        compress_module compress_581 (
                                            .x(u[2][69]),
                                            .d(10),
                                            .result(com_out[2][69])
                                        );
                                        
                                        compress_module compress_582 (
                                            .x(u[2][70]),
                                            .d(10),
                                            .result(com_out[2][70])
                                        );
                                        
                                        compress_module compress_583 (
                                            .x(u[2][71]),
                                            .d(10),
                                            .result(com_out[2][71])
                                        );
                                        
                                        compress_module compress_584 (
                                            .x(u[2][72]),
                                            .d(10),
                                            .result(com_out[2][72])
                                        );
                                        
                                        compress_module compress_585 (
                                            .x(u[2][73]),
                                            .d(10),
                                            .result(com_out[2][73])
                                        );
                                        
                                        compress_module compress_586 (
                                            .x(u[2][74]),
                                            .d(10),
                                            .result(com_out[2][74])
                                        );
                                        
                                        compress_module compress_587 (
                                            .x(u[2][75]),
                                            .d(10),
                                            .result(com_out[2][75])
                                        );
                                        
                                        compress_module compress_588 (
                                            .x(u[2][76]),
                                            .d(10),
                                            .result(com_out[2][76])
                                        );
                                        
                                        compress_module compress_589 (
                                            .x(u[2][77]),
                                            .d(10),
                                            .result(com_out[2][77])
                                        );
                                        
                                        compress_module compress_590 (
                                            .x(u[2][78]),
                                            .d(10),
                                            .result(com_out[2][78])
                                        );
                                        
                                        compress_module compress_591 (
                                            .x(u[2][79]),
                                            .d(10),
                                            .result(com_out[2][79])
                                        );
                                        
                                        compress_module compress_592 (
                                            .x(u[2][80]),
                                            .d(10),
                                            .result(com_out[2][80])
                                        );
                                        
                                        compress_module compress_593 (
                                            .x(u[2][81]),
                                            .d(10),
                                            .result(com_out[2][81])
                                        );
                                        
                                        compress_module compress_594 (
                                            .x(u[2][82]),
                                            .d(10),
                                            .result(com_out[2][82])
                                        );
                                        
                                        compress_module compress_595 (
                                            .x(u[2][83]),
                                            .d(10),
                                            .result(com_out[2][83])
                                        );
                                        
                                        compress_module compress_596 (
                                            .x(u[2][84]),
                                            .d(10),
                                            .result(com_out[2][84])
                                        );
                                        
                                        compress_module compress_597 (
                                            .x(u[2][85]),
                                            .d(10),
                                            .result(com_out[2][85])
                                        );
                                        
                                        compress_module compress_598 (
                                            .x(u[2][86]),
                                            .d(10),
                                            .result(com_out[2][86])
                                        );
                                        
                                        compress_module compress_599 (
                                            .x(u[2][87]),
                                            .d(10),
                                            .result(com_out[2][87])
                                        );
                                        
                                        compress_module compress_600 (
                                            .x(u[2][88]),
                                            .d(10),
                                            .result(com_out[2][88])
                                        );
                                        
                                        compress_module compress_601 (
                                            .x(u[2][89]),
                                            .d(10),
                                            .result(com_out[2][89])
                                        );
                                        
                                        compress_module compress_602 (
                                            .x(u[2][90]),
                                            .d(10),
                                            .result(com_out[2][90])
                                        );
                                        
                                        compress_module compress_603 (
                                            .x(u[2][91]),
                                            .d(10),
                                            .result(com_out[2][91])
                                        );
                                        
                                        compress_module compress_604 (
                                            .x(u[2][92]),
                                            .d(10),
                                            .result(com_out[2][92])
                                        );
                                        
                                        compress_module compress_605 (
                                            .x(u[2][93]),
                                            .d(10),
                                            .result(com_out[2][93])
                                        );
                                        
                                        compress_module compress_606 (
                                            .x(u[2][94]),
                                            .d(10),
                                            .result(com_out[2][94])
                                        );
                                        
                                        compress_module compress_607 (
                                            .x(u[2][95]),
                                            .d(10),
                                            .result(com_out[2][95])
                                        );
                                        
                                        compress_module compress_608 (
                                            .x(u[2][96]),
                                            .d(10),
                                            .result(com_out[2][96])
                                        );
                                        
                                        compress_module compress_609 (
                                            .x(u[2][97]),
                                            .d(10),
                                            .result(com_out[2][97])
                                        );
                                        
                                        compress_module compress_610 (
                                            .x(u[2][98]),
                                            .d(10),
                                            .result(com_out[2][98])
                                        );
                                        
                                        compress_module compress_611 (
                                            .x(u[2][99]),
                                            .d(10),
                                            .result(com_out[2][99])
                                        );
                                        
                                        compress_module compress_612 (
                                            .x(u[2][100]),
                                            .d(10),
                                            .result(com_out[2][100])
                                        );
                                        
                                        compress_module compress_613 (
                                            .x(u[2][101]),
                                            .d(10),
                                            .result(com_out[2][101])
                                        );
                                        
                                        compress_module compress_614 (
                                            .x(u[2][102]),
                                            .d(10),
                                            .result(com_out[2][102])
                                        );
                                        
                                        compress_module compress_615 (
                                            .x(u[2][103]),
                                            .d(10),
                                            .result(com_out[2][103])
                                        );
                                        
                                        compress_module compress_616 (
                                            .x(u[2][104]),
                                            .d(10),
                                            .result(com_out[2][104])
                                        );
                                        
                                        compress_module compress_617 (
                                            .x(u[2][105]),
                                            .d(10),
                                            .result(com_out[2][105])
                                        );
                                        
                                        compress_module compress_618 (
                                            .x(u[2][106]),
                                            .d(10),
                                            .result(com_out[2][106])
                                        );
                                        
                                        compress_module compress_619 (
                                            .x(u[2][107]),
                                            .d(10),
                                            .result(com_out[2][107])
                                        );
                                        
                                        compress_module compress_620 (
                                            .x(u[2][108]),
                                            .d(10),
                                            .result(com_out[2][108])
                                        );
                                        
                                        compress_module compress_621 (
                                            .x(u[2][109]),
                                            .d(10),
                                            .result(com_out[2][109])
                                        );
                                        
                                        compress_module compress_622 (
                                            .x(u[2][110]),
                                            .d(10),
                                            .result(com_out[2][110])
                                        );
                                        
                                        compress_module compress_623 (
                                            .x(u[2][111]),
                                            .d(10),
                                            .result(com_out[2][111])
                                        );
                                        
                                        compress_module compress_624 (
                                            .x(u[2][112]),
                                            .d(10),
                                            .result(com_out[2][112])
                                        );
                                        
                                        compress_module compress_625 (
                                            .x(u[2][113]),
                                            .d(10),
                                            .result(com_out[2][113])
                                        );
                                        
                                        compress_module compress_626 (
                                            .x(u[2][114]),
                                            .d(10),
                                            .result(com_out[2][114])
                                        );
                                        
                                        compress_module compress_627 (
                                            .x(u[2][115]),
                                            .d(10),
                                            .result(com_out[2][115])
                                        );
                                        
                                        compress_module compress_628 (
                                            .x(u[2][116]),
                                            .d(10),
                                            .result(com_out[2][116])
                                        );
                                        
                                        compress_module compress_629 (
                                            .x(u[2][117]),
                                            .d(10),
                                            .result(com_out[2][117])
                                        );
                                        
                                        compress_module compress_630 (
                                            .x(u[2][118]),
                                            .d(10),
                                            .result(com_out[2][118])
                                        );
                                        
                                        compress_module compress_631 (
                                            .x(u[2][119]),
                                            .d(10),
                                            .result(com_out[2][119])
                                        );
                                        
                                        compress_module compress_632 (
                                            .x(u[2][120]),
                                            .d(10),
                                            .result(com_out[2][120])
                                        );
                                        
                                        compress_module compress_633 (
                                            .x(u[2][121]),
                                            .d(10),
                                            .result(com_out[2][121])
                                        );
                                        
                                        compress_module compress_634 (
                                            .x(u[2][122]),
                                            .d(10),
                                            .result(com_out[2][122])
                                        );
                                        
                                        compress_module compress_635 (
                                            .x(u[2][123]),
                                            .d(10),
                                            .result(com_out[2][123])
                                        );
                                        
                                        compress_module compress_636 (
                                            .x(u[2][124]),
                                            .d(10),
                                            .result(com_out[2][124])
                                        );
                                        
                                        compress_module compress_637 (
                                            .x(u[2][125]),
                                            .d(10),
                                            .result(com_out[2][125])
                                        );
                                        
                                        compress_module compress_638 (
                                            .x(u[2][126]),
                                            .d(10),
                                            .result(com_out[2][126])
                                        );
                                        
                                        compress_module compress_639 (
                                            .x(u[2][127]),
                                            .d(10),
                                            .result(com_out[2][127])
                                        );
                                        
                                        compress_module compress_640 (
                                            .x(u[2][128]),
                                            .d(10),
                                            .result(com_out[2][128])
                                        );
                                        
                                        compress_module compress_641 (
                                            .x(u[2][129]),
                                            .d(10),
                                            .result(com_out[2][129])
                                        );
                                        
                                        compress_module compress_642 (
                                            .x(u[2][130]),
                                            .d(10),
                                            .result(com_out[2][130])
                                        );
                                        
                                        compress_module compress_643 (
                                            .x(u[2][131]),
                                            .d(10),
                                            .result(com_out[2][131])
                                        );
                                        
                                        compress_module compress_644 (
                                            .x(u[2][132]),
                                            .d(10),
                                            .result(com_out[2][132])
                                        );
                                        
                                        compress_module compress_645 (
                                            .x(u[2][133]),
                                            .d(10),
                                            .result(com_out[2][133])
                                        );
                                        
                                        compress_module compress_646 (
                                            .x(u[2][134]),
                                            .d(10),
                                            .result(com_out[2][134])
                                        );
                                        
                                        compress_module compress_647 (
                                            .x(u[2][135]),
                                            .d(10),
                                            .result(com_out[2][135])
                                        );
                                        
                                        compress_module compress_648 (
                                            .x(u[2][136]),
                                            .d(10),
                                            .result(com_out[2][136])
                                        );
                                        
                                        compress_module compress_649 (
                                            .x(u[2][137]),
                                            .d(10),
                                            .result(com_out[2][137])
                                        );
                                        
                                        compress_module compress_650 (
                                            .x(u[2][138]),
                                            .d(10),
                                            .result(com_out[2][138])
                                        );
                                        
                                        compress_module compress_651 (
                                            .x(u[2][139]),
                                            .d(10),
                                            .result(com_out[2][139])
                                        );
                                        
                                        compress_module compress_652 (
                                            .x(u[2][140]),
                                            .d(10),
                                            .result(com_out[2][140])
                                        );
                                        
                                        compress_module compress_653 (
                                            .x(u[2][141]),
                                            .d(10),
                                            .result(com_out[2][141])
                                        );
                                        
                                        compress_module compress_654 (
                                            .x(u[2][142]),
                                            .d(10),
                                            .result(com_out[2][142])
                                        );
                                        
                                        compress_module compress_655 (
                                            .x(u[2][143]),
                                            .d(10),
                                            .result(com_out[2][143])
                                        );
                                        
                                        compress_module compress_656 (
                                            .x(u[2][144]),
                                            .d(10),
                                            .result(com_out[2][144])
                                        );
                                        
                                        compress_module compress_657 (
                                            .x(u[2][145]),
                                            .d(10),
                                            .result(com_out[2][145])
                                        );
                                        
                                        compress_module compress_658 (
                                            .x(u[2][146]),
                                            .d(10),
                                            .result(com_out[2][146])
                                        );
                                        
                                        compress_module compress_659 (
                                            .x(u[2][147]),
                                            .d(10),
                                            .result(com_out[2][147])
                                        );
                                        
                                        compress_module compress_660 (
                                            .x(u[2][148]),
                                            .d(10),
                                            .result(com_out[2][148])
                                        );
                                        
                                        compress_module compress_661 (
                                            .x(u[2][149]),
                                            .d(10),
                                            .result(com_out[2][149])
                                        );
                                        
                                        compress_module compress_662 (
                                            .x(u[2][150]),
                                            .d(10),
                                            .result(com_out[2][150])
                                        );
                                        
                                        compress_module compress_663 (
                                            .x(u[2][151]),
                                            .d(10),
                                            .result(com_out[2][151])
                                        );
                                        
                                        compress_module compress_664 (
                                            .x(u[2][152]),
                                            .d(10),
                                            .result(com_out[2][152])
                                        );
                                        
                                        compress_module compress_665 (
                                            .x(u[2][153]),
                                            .d(10),
                                            .result(com_out[2][153])
                                        );
                                        
                                        compress_module compress_666 (
                                            .x(u[2][154]),
                                            .d(10),
                                            .result(com_out[2][154])
                                        );
                                        
                                        compress_module compress_667 (
                                            .x(u[2][155]),
                                            .d(10),
                                            .result(com_out[2][155])
                                        );
                                        
                                        compress_module compress_668 (
                                            .x(u[2][156]),
                                            .d(10),
                                            .result(com_out[2][156])
                                        );
                                        
                                        compress_module compress_669 (
                                            .x(u[2][157]),
                                            .d(10),
                                            .result(com_out[2][157])
                                        );
                                        
                                        compress_module compress_670 (
                                            .x(u[2][158]),
                                            .d(10),
                                            .result(com_out[2][158])
                                        );
                                        
                                        compress_module compress_671 (
                                            .x(u[2][159]),
                                            .d(10),
                                            .result(com_out[2][159])
                                        );
                                        
                                        compress_module compress_672 (
                                            .x(u[2][160]),
                                            .d(10),
                                            .result(com_out[2][160])
                                        );
                                        
                                        compress_module compress_673 (
                                            .x(u[2][161]),
                                            .d(10),
                                            .result(com_out[2][161])
                                        );
                                        
                                        compress_module compress_674 (
                                            .x(u[2][162]),
                                            .d(10),
                                            .result(com_out[2][162])
                                        );
                                        
                                        compress_module compress_675 (
                                            .x(u[2][163]),
                                            .d(10),
                                            .result(com_out[2][163])
                                        );
                                        
                                        compress_module compress_676 (
                                            .x(u[2][164]),
                                            .d(10),
                                            .result(com_out[2][164])
                                        );
                                        
                                        compress_module compress_677 (
                                            .x(u[2][165]),
                                            .d(10),
                                            .result(com_out[2][165])
                                        );
                                        
                                        compress_module compress_678 (
                                            .x(u[2][166]),
                                            .d(10),
                                            .result(com_out[2][166])
                                        );
                                        
                                        compress_module compress_679 (
                                            .x(u[2][167]),
                                            .d(10),
                                            .result(com_out[2][167])
                                        );
                                        
                                        compress_module compress_680 (
                                            .x(u[2][168]),
                                            .d(10),
                                            .result(com_out[2][168])
                                        );
                                        
                                        compress_module compress_681 (
                                            .x(u[2][169]),
                                            .d(10),
                                            .result(com_out[2][169])
                                        );
                                        
                                        compress_module compress_682 (
                                            .x(u[2][170]),
                                            .d(10),
                                            .result(com_out[2][170])
                                        );
                                        
                                        compress_module compress_683 (
                                            .x(u[2][171]),
                                            .d(10),
                                            .result(com_out[2][171])
                                        );
                                        
                                        compress_module compress_684 (
                                            .x(u[2][172]),
                                            .d(10),
                                            .result(com_out[2][172])
                                        );
                                        
                                        compress_module compress_685 (
                                            .x(u[2][173]),
                                            .d(10),
                                            .result(com_out[2][173])
                                        );
                                        
                                        compress_module compress_686 (
                                            .x(u[2][174]),
                                            .d(10),
                                            .result(com_out[2][174])
                                        );
                                        
                                        compress_module compress_687 (
                                            .x(u[2][175]),
                                            .d(10),
                                            .result(com_out[2][175])
                                        );
                                        
                                        compress_module compress_688 (
                                            .x(u[2][176]),
                                            .d(10),
                                            .result(com_out[2][176])
                                        );
                                        
                                        compress_module compress_689 (
                                            .x(u[2][177]),
                                            .d(10),
                                            .result(com_out[2][177])
                                        );
                                        
                                        compress_module compress_690 (
                                            .x(u[2][178]),
                                            .d(10),
                                            .result(com_out[2][178])
                                        );
                                        
                                        compress_module compress_691 (
                                            .x(u[2][179]),
                                            .d(10),
                                            .result(com_out[2][179])
                                        );
                                        
                                        compress_module compress_692 (
                                            .x(u[2][180]),
                                            .d(10),
                                            .result(com_out[2][180])
                                        );
                                        
                                        compress_module compress_693 (
                                            .x(u[2][181]),
                                            .d(10),
                                            .result(com_out[2][181])
                                        );
                                        
                                        compress_module compress_694 (
                                            .x(u[2][182]),
                                            .d(10),
                                            .result(com_out[2][182])
                                        );
                                        
                                        compress_module compress_695 (
                                            .x(u[2][183]),
                                            .d(10),
                                            .result(com_out[2][183])
                                        );
                                        
                                        compress_module compress_696 (
                                            .x(u[2][184]),
                                            .d(10),
                                            .result(com_out[2][184])
                                        );
                                        
                                        compress_module compress_697 (
                                            .x(u[2][185]),
                                            .d(10),
                                            .result(com_out[2][185])
                                        );
                                        
                                        compress_module compress_698 (
                                            .x(u[2][186]),
                                            .d(10),
                                            .result(com_out[2][186])
                                        );
                                        
                                        compress_module compress_699 (
                                            .x(u[2][187]),
                                            .d(10),
                                            .result(com_out[2][187])
                                        );
                                        
                                        compress_module compress_700 (
                                            .x(u[2][188]),
                                            .d(10),
                                            .result(com_out[2][188])
                                        );
                                        
                                        compress_module compress_701 (
                                            .x(u[2][189]),
                                            .d(10),
                                            .result(com_out[2][189])
                                        );
                                        
                                        compress_module compress_702 (
                                            .x(u[2][190]),
                                            .d(10),
                                            .result(com_out[2][190])
                                        );
                                        
                                        compress_module compress_703 (
                                            .x(u[2][191]),
                                            .d(10),
                                            .result(com_out[2][191])
                                        );
                                        
                                        compress_module compress_704 (
                                            .x(u[2][192]),
                                            .d(10),
                                            .result(com_out[2][192])
                                        );
                                        
                                        compress_module compress_705 (
                                            .x(u[2][193]),
                                            .d(10),
                                            .result(com_out[2][193])
                                        );
                                        
                                        compress_module compress_706 (
                                            .x(u[2][194]),
                                            .d(10),
                                            .result(com_out[2][194])
                                        );
                                        
                                        compress_module compress_707 (
                                            .x(u[2][195]),
                                            .d(10),
                                            .result(com_out[2][195])
                                        );
                                        
                                        compress_module compress_708 (
                                            .x(u[2][196]),
                                            .d(10),
                                            .result(com_out[2][196])
                                        );
                                        
                                        compress_module compress_709 (
                                            .x(u[2][197]),
                                            .d(10),
                                            .result(com_out[2][197])
                                        );
                                        
                                        compress_module compress_710 (
                                            .x(u[2][198]),
                                            .d(10),
                                            .result(com_out[2][198])
                                        );
                                        
                                        compress_module compress_711 (
                                            .x(u[2][199]),
                                            .d(10),
                                            .result(com_out[2][199])
                                        );
                                        
                                        compress_module compress_712 (
                                            .x(u[2][200]),
                                            .d(10),
                                            .result(com_out[2][200])
                                        );
                                        
                                        compress_module compress_713 (
                                            .x(u[2][201]),
                                            .d(10),
                                            .result(com_out[2][201])
                                        );
                                        
                                        compress_module compress_714 (
                                            .x(u[2][202]),
                                            .d(10),
                                            .result(com_out[2][202])
                                        );
                                        
                                        compress_module compress_715 (
                                            .x(u[2][203]),
                                            .d(10),
                                            .result(com_out[2][203])
                                        );
                                        
                                        compress_module compress_716 (
                                            .x(u[2][204]),
                                            .d(10),
                                            .result(com_out[2][204])
                                        );
                                        
                                        compress_module compress_717 (
                                            .x(u[2][205]),
                                            .d(10),
                                            .result(com_out[2][205])
                                        );
                                        
                                        compress_module compress_718 (
                                            .x(u[2][206]),
                                            .d(10),
                                            .result(com_out[2][206])
                                        );
                                        
                                        compress_module compress_719 (
                                            .x(u[2][207]),
                                            .d(10),
                                            .result(com_out[2][207])
                                        );
                                        
                                        compress_module compress_720 (
                                            .x(u[2][208]),
                                            .d(10),
                                            .result(com_out[2][208])
                                        );
                                        
                                        compress_module compress_721 (
                                            .x(u[2][209]),
                                            .d(10),
                                            .result(com_out[2][209])
                                        );
                                        
                                        compress_module compress_722 (
                                            .x(u[2][210]),
                                            .d(10),
                                            .result(com_out[2][210])
                                        );
                                        
                                        compress_module compress_723 (
                                            .x(u[2][211]),
                                            .d(10),
                                            .result(com_out[2][211])
                                        );
                                        
                                        compress_module compress_724 (
                                            .x(u[2][212]),
                                            .d(10),
                                            .result(com_out[2][212])
                                        );
                                        
                                        compress_module compress_725 (
                                            .x(u[2][213]),
                                            .d(10),
                                            .result(com_out[2][213])
                                        );
                                        
                                        compress_module compress_726 (
                                            .x(u[2][214]),
                                            .d(10),
                                            .result(com_out[2][214])
                                        );
                                        
                                        compress_module compress_727 (
                                            .x(u[2][215]),
                                            .d(10),
                                            .result(com_out[2][215])
                                        );
                                        
                                        compress_module compress_728 (
                                            .x(u[2][216]),
                                            .d(10),
                                            .result(com_out[2][216])
                                        );
                                        
                                        compress_module compress_729 (
                                            .x(u[2][217]),
                                            .d(10),
                                            .result(com_out[2][217])
                                        );
                                        
                                        compress_module compress_730 (
                                            .x(u[2][218]),
                                            .d(10),
                                            .result(com_out[2][218])
                                        );
                                        
                                        compress_module compress_731 (
                                            .x(u[2][219]),
                                            .d(10),
                                            .result(com_out[2][219])
                                        );
                                        
                                        compress_module compress_732 (
                                            .x(u[2][220]),
                                            .d(10),
                                            .result(com_out[2][220])
                                        );
                                        
                                        compress_module compress_733 (
                                            .x(u[2][221]),
                                            .d(10),
                                            .result(com_out[2][221])
                                        );
                                        
                                        compress_module compress_734 (
                                            .x(u[2][222]),
                                            .d(10),
                                            .result(com_out[2][222])
                                        );
                                        
                                        compress_module compress_735 (
                                            .x(u[2][223]),
                                            .d(10),
                                            .result(com_out[2][223])
                                        );
                                        
                                        compress_module compress_736 (
                                            .x(u[2][224]),
                                            .d(10),
                                            .result(com_out[2][224])
                                        );
                                        
                                        compress_module compress_737 (
                                            .x(u[2][225]),
                                            .d(10),
                                            .result(com_out[2][225])
                                        );
                                        
                                        compress_module compress_738 (
                                            .x(u[2][226]),
                                            .d(10),
                                            .result(com_out[2][226])
                                        );
                                        
                                        compress_module compress_739 (
                                            .x(u[2][227]),
                                            .d(10),
                                            .result(com_out[2][227])
                                        );
                                        
                                        compress_module compress_740 (
                                            .x(u[2][228]),
                                            .d(10),
                                            .result(com_out[2][228])
                                        );
                                        
                                        compress_module compress_741 (
                                            .x(u[2][229]),
                                            .d(10),
                                            .result(com_out[2][229])
                                        );
                                        
                                        compress_module compress_742 (
                                            .x(u[2][230]),
                                            .d(10),
                                            .result(com_out[2][230])
                                        );
                                        
                                        compress_module compress_743 (
                                            .x(u[2][231]),
                                            .d(10),
                                            .result(com_out[2][231])
                                        );
                                        
                                        compress_module compress_744 (
                                            .x(u[2][232]),
                                            .d(10),
                                            .result(com_out[2][232])
                                        );
                                        
                                        compress_module compress_745 (
                                            .x(u[2][233]),
                                            .d(10),
                                            .result(com_out[2][233])
                                        );
                                        
                                        compress_module compress_746 (
                                            .x(u[2][234]),
                                            .d(10),
                                            .result(com_out[2][234])
                                        );
                                        
                                        compress_module compress_747 (
                                            .x(u[2][235]),
                                            .d(10),
                                            .result(com_out[2][235])
                                        );
                                        
                                        compress_module compress_748 (
                                            .x(u[2][236]),
                                            .d(10),
                                            .result(com_out[2][236])
                                        );
                                        
                                        compress_module compress_749 (
                                            .x(u[2][237]),
                                            .d(10),
                                            .result(com_out[2][237])
                                        );
                                        
                                        compress_module compress_750 (
                                            .x(u[2][238]),
                                            .d(10),
                                            .result(com_out[2][238])
                                        );
                                        
                                        compress_module compress_751 (
                                            .x(u[2][239]),
                                            .d(10),
                                            .result(com_out[2][239])
                                        );
                                        
                                        compress_module compress_752 (
                                            .x(u[2][240]),
                                            .d(10),
                                            .result(com_out[2][240])
                                        );
                                        
                                        compress_module compress_753 (
                                            .x(u[2][241]),
                                            .d(10),
                                            .result(com_out[2][241])
                                        );
                                        
                                        compress_module compress_754 (
                                            .x(u[2][242]),
                                            .d(10),
                                            .result(com_out[2][242])
                                        );
                                        
                                        compress_module compress_755 (
                                            .x(u[2][243]),
                                            .d(10),
                                            .result(com_out[2][243])
                                        );
                                        
                                        compress_module compress_756 (
                                            .x(u[2][244]),
                                            .d(10),
                                            .result(com_out[2][244])
                                        );
                                        
                                        compress_module compress_757 (
                                            .x(u[2][245]),
                                            .d(10),
                                            .result(com_out[2][245])
                                        );
                                        
                                        compress_module compress_758 (
                                            .x(u[2][246]),
                                            .d(10),
                                            .result(com_out[2][246])
                                        );
                                        
                                        compress_module compress_759 (
                                            .x(u[2][247]),
                                            .d(10),
                                            .result(com_out[2][247])
                                        );
                                        
                                        compress_module compress_760 (
                                            .x(u[2][248]),
                                            .d(10),
                                            .result(com_out[2][248])
                                        );
                                        
                                        compress_module compress_761 (
                                            .x(u[2][249]),
                                            .d(10),
                                            .result(com_out[2][249])
                                        );
                                        
                                        compress_module compress_762 (
                                            .x(u[2][250]),
                                            .d(10),
                                            .result(com_out[2][250])
                                        );
                                        
                                        compress_module compress_763 (
                                            .x(u[2][251]),
                                            .d(10),
                                            .result(com_out[2][251])
                                        );
                                        
                                        compress_module compress_764 (
                                            .x(u[2][252]),
                                            .d(10),
                                            .result(com_out[2][252])
                                        );
                                        
                                        compress_module compress_765 (
                                            .x(u[2][253]),
                                            .d(10),
                                            .result(com_out[2][253])
                                        );
                                        
                                        compress_module compress_766 (
                                            .x(u[2][254]),
                                            .d(10),
                                            .result(com_out[2][254])
                                        );
                                        
                                        compress_module compress_767 (
                                            .x(u[2][255]),
                                            .d(10),
                                            .result(com_out[2][255])
                                        );
                                       compress_module comp_v_0 (
                                            .x(v[0]),
                                            .d(4),
                                            .result(comp_v[0])
                                        );
                                        
                                        compress_module comp_v_1 (
                                            .x(v[1]),
                                            .d(4),
                                            .result(comp_v[1])
                                        );
                                        
                                        compress_module comp_v_2 (
                                            .x(v[2]),
                                            .d(4),
                                            .result(comp_v[2])
                                        );
                                        
                                        compress_module comp_v_3 (
                                            .x(v[3]),
                                            .d(4),
                                            .result(comp_v[3])
                                        );
                                        
                                        compress_module comp_v_4 (
                                            .x(v[4]),
                                            .d(4),
                                            .result(comp_v[4])
                                        );
                                        
                                        compress_module comp_v_5 (
                                            .x(v[5]),
                                            .d(4),
                                            .result(comp_v[5])
                                        );
                                        
                                        compress_module comp_v_6 (
                                            .x(v[6]),
                                            .d(4),
                                            .result(comp_v[6])
                                        );
                                        
                                        compress_module comp_v_7 (
                                            .x(v[7]),
                                            .d(4),
                                            .result(comp_v[7])
                                        );
                                        
                                        compress_module comp_v_8 (
                                            .x(v[8]),
                                            .d(4),
                                            .result(comp_v[8])
                                        );
                                        
                                        compress_module comp_v_9 (
                                            .x(v[9]),
                                            .d(4),
                                            .result(comp_v[9])
                                        );
                                        
                                        compress_module comp_v_10 (
                                            .x(v[10]),
                                            .d(4),
                                            .result(comp_v[10])
                                        );
                                        
                                        compress_module comp_v_11 (
                                            .x(v[11]),
                                            .d(4),
                                            .result(comp_v[11])
                                        );
                                        
                                        compress_module comp_v_12 (
                                            .x(v[12]),
                                            .d(4),
                                            .result(comp_v[12])
                                        );
                                        
                                        compress_module comp_v_13 (
                                            .x(v[13]),
                                            .d(4),
                                            .result(comp_v[13])
                                        );
                                        
                                        compress_module comp_v_14 (
                                            .x(v[14]),
                                            .d(4),
                                            .result(comp_v[14])
                                        );
                                        
                                        compress_module comp_v_15 (
                                            .x(v[15]),
                                            .d(4),
                                            .result(comp_v[15])
                                        );
                                        
                                        compress_module comp_v_16 (
                                            .x(v[16]),
                                            .d(4),
                                            .result(comp_v[16])
                                        );
                                        
                                        compress_module comp_v_17 (
                                            .x(v[17]),
                                            .d(4),
                                            .result(comp_v[17])
                                        );
                                        
                                        compress_module comp_v_18 (
                                            .x(v[18]),
                                            .d(4),
                                            .result(comp_v[18])
                                        );
                                        
                                        compress_module comp_v_19 (
                                            .x(v[19]),
                                            .d(4),
                                            .result(comp_v[19])
                                        );
                                        
                                        compress_module comp_v_20 (
                                            .x(v[20]),
                                            .d(4),
                                            .result(comp_v[20])
                                        );
                                        
                                        compress_module comp_v_21 (
                                            .x(v[21]),
                                            .d(4),
                                            .result(comp_v[21])
                                        );
                                        
                                        compress_module comp_v_22 (
                                            .x(v[22]),
                                            .d(4),
                                            .result(comp_v[22])
                                        );
                                        
                                        compress_module comp_v_23 (
                                            .x(v[23]),
                                            .d(4),
                                            .result(comp_v[23])
                                        );
                                        
                                        compress_module comp_v_24 (
                                            .x(v[24]),
                                            .d(4),
                                            .result(comp_v[24])
                                        );
                                        
                                        compress_module comp_v_25 (
                                            .x(v[25]),
                                            .d(4),
                                            .result(comp_v[25])
                                        );
                                        
                                        compress_module comp_v_26 (
                                            .x(v[26]),
                                            .d(4),
                                            .result(comp_v[26])
                                        );
                                        
                                        compress_module comp_v_27 (
                                            .x(v[27]),
                                            .d(4),
                                            .result(comp_v[27])
                                        );
                                        
                                        compress_module comp_v_28 (
                                            .x(v[28]),
                                            .d(4),
                                            .result(comp_v[28])
                                        );
                                        
                                        compress_module comp_v_29 (
                                            .x(v[29]),
                                            .d(4),
                                            .result(comp_v[29])
                                        );
                                        
                                        compress_module comp_v_30 (
                                            .x(v[30]),
                                            .d(4),
                                            .result(comp_v[30])
                                        );
                                        
                                        compress_module comp_v_31 (
                                            .x(v[31]),
                                            .d(4),
                                            .result(comp_v[31])
                                        );
                                        
                                        compress_module comp_v_32 (
                                            .x(v[32]),
                                            .d(4),
                                            .result(comp_v[32])
                                        );
                                        
                                        compress_module comp_v_33 (
                                            .x(v[33]),
                                            .d(4),
                                            .result(comp_v[33])
                                        );
                                        
                                        compress_module comp_v_34 (
                                            .x(v[34]),
                                            .d(4),
                                            .result(comp_v[34])
                                        );
                                        
                                        compress_module comp_v_35 (
                                            .x(v[35]),
                                            .d(4),
                                            .result(comp_v[35])
                                        );
                                        
                                        compress_module comp_v_36 (
                                            .x(v[36]),
                                            .d(4),
                                            .result(comp_v[36])
                                        );
                                        
                                        compress_module comp_v_37 (
                                            .x(v[37]),
                                            .d(4),
                                            .result(comp_v[37])
                                        );
                                        
                                        compress_module comp_v_38 (
                                            .x(v[38]),
                                            .d(4),
                                            .result(comp_v[38])
                                        );
                                        
                                        compress_module comp_v_39 (
                                            .x(v[39]),
                                            .d(4),
                                            .result(comp_v[39])
                                        );
                                        
                                        compress_module comp_v_40 (
                                            .x(v[40]),
                                            .d(4),
                                            .result(comp_v[40])
                                        );
                                        
                                        compress_module comp_v_41 (
                                            .x(v[41]),
                                            .d(4),
                                            .result(comp_v[41])
                                        );
                                        
                                        compress_module comp_v_42 (
                                            .x(v[42]),
                                            .d(4),
                                            .result(comp_v[42])
                                        );
                                        
                                        compress_module comp_v_43 (
                                            .x(v[43]),
                                            .d(4),
                                            .result(comp_v[43])
                                        );
                                        
                                        compress_module comp_v_44 (
                                            .x(v[44]),
                                            .d(4),
                                            .result(comp_v[44])
                                        );
                                        
                                        compress_module comp_v_45 (
                                            .x(v[45]),
                                            .d(4),
                                            .result(comp_v[45])
                                        );
                                        
                                        compress_module comp_v_46 (
                                            .x(v[46]),
                                            .d(4),
                                            .result(comp_v[46])
                                        );
                                        
                                        compress_module comp_v_47 (
                                            .x(v[47]),
                                            .d(4),
                                            .result(comp_v[47])
                                        );
                                        
                                        compress_module comp_v_48 (
                                            .x(v[48]),
                                            .d(4),
                                            .result(comp_v[48])
                                        );
                                        
                                        compress_module comp_v_49 (
                                            .x(v[49]),
                                            .d(4),
                                            .result(comp_v[49])
                                        );
                                        
                                        compress_module comp_v_50 (
                                            .x(v[50]),
                                            .d(4),
                                            .result(comp_v[50])
                                        );
                                        
                                        compress_module comp_v_51 (
                                            .x(v[51]),
                                            .d(4),
                                            .result(comp_v[51])
                                        );
                                        
                                        compress_module comp_v_52 (
                                            .x(v[52]),
                                            .d(4),
                                            .result(comp_v[52])
                                        );
                                        
                                        compress_module comp_v_53 (
                                            .x(v[53]),
                                            .d(4),
                                            .result(comp_v[53])
                                        );
                                        
                                        compress_module comp_v_54 (
                                            .x(v[54]),
                                            .d(4),
                                            .result(comp_v[54])
                                        );
                                        
                                        compress_module comp_v_55 (
                                            .x(v[55]),
                                            .d(4),
                                            .result(comp_v[55])
                                        );
                                        
                                        compress_module comp_v_56 (
                                            .x(v[56]),
                                            .d(4),
                                            .result(comp_v[56])
                                        );
                                        
                                        compress_module comp_v_57 (
                                            .x(v[57]),
                                            .d(4),
                                            .result(comp_v[57])
                                        );
                                        
                                        compress_module comp_v_58 (
                                            .x(v[58]),
                                            .d(4),
                                            .result(comp_v[58])
                                        );
                                        
                                        compress_module comp_v_59 (
                                            .x(v[59]),
                                            .d(4),
                                            .result(comp_v[59])
                                        );
                                        
                                        compress_module comp_v_60 (
                                            .x(v[60]),
                                            .d(4),
                                            .result(comp_v[60])
                                        );
                                        
                                        compress_module comp_v_61 (
                                            .x(v[61]),
                                            .d(4),
                                            .result(comp_v[61])
                                        );
                                        
                                        compress_module comp_v_62 (
                                            .x(v[62]),
                                            .d(4),
                                            .result(comp_v[62])
                                        );
                                        
                                        compress_module comp_v_63 (
                                            .x(v[63]),
                                            .d(4),
                                            .result(comp_v[63])
                                        );
                                        
                                        compress_module comp_v_64 (
                                            .x(v[64]),
                                            .d(4),
                                            .result(comp_v[64])
                                        );
                                        
                                        compress_module comp_v_65 (
                                            .x(v[65]),
                                            .d(4),
                                            .result(comp_v[65])
                                        );
                                        
                                        compress_module comp_v_66 (
                                            .x(v[66]),
                                            .d(4),
                                            .result(comp_v[66])
                                        );
                                        
                                        compress_module comp_v_67 (
                                            .x(v[67]),
                                            .d(4),
                                            .result(comp_v[67])
                                        );
                                        
                                        compress_module comp_v_68 (
                                            .x(v[68]),
                                            .d(4),
                                            .result(comp_v[68])
                                        );
                                        
                                        compress_module comp_v_69 (
                                            .x(v[69]),
                                            .d(4),
                                            .result(comp_v[69])
                                        );
                                        
                                        compress_module comp_v_70 (
                                            .x(v[70]),
                                            .d(4),
                                            .result(comp_v[70])
                                        );
                                        
                                        compress_module comp_v_71 (
                                            .x(v[71]),
                                            .d(4),
                                            .result(comp_v[71])
                                        );
                                        
                                        compress_module comp_v_72 (
                                            .x(v[72]),
                                            .d(4),
                                            .result(comp_v[72])
                                        );
                                        
                                        compress_module comp_v_73 (
                                            .x(v[73]),
                                            .d(4),
                                            .result(comp_v[73])
                                        );
                                        
                                        compress_module comp_v_74 (
                                            .x(v[74]),
                                            .d(4),
                                            .result(comp_v[74])
                                        );
                                        
                                        compress_module comp_v_75 (
                                            .x(v[75]),
                                            .d(4),
                                            .result(comp_v[75])
                                        );
                                        
                                        compress_module comp_v_76 (
                                            .x(v[76]),
                                            .d(4),
                                            .result(comp_v[76])
                                        );
                                        
                                        compress_module comp_v_77 (
                                            .x(v[77]),
                                            .d(4),
                                            .result(comp_v[77])
                                        );
                                        
                                        compress_module comp_v_78 (
                                            .x(v[78]),
                                            .d(4),
                                            .result(comp_v[78])
                                        );
                                        
                                        compress_module comp_v_79 (
                                            .x(v[79]),
                                            .d(4),
                                            .result(comp_v[79])
                                        );
                                        
                                        compress_module comp_v_80 (
                                            .x(v[80]),
                                            .d(4),
                                            .result(comp_v[80])
                                        );
                                        
                                        compress_module comp_v_81 (
                                            .x(v[81]),
                                            .d(4),
                                            .result(comp_v[81])
                                        );
                                        
                                        compress_module comp_v_82 (
                                            .x(v[82]),
                                            .d(4),
                                            .result(comp_v[82])
                                        );
                                        
                                        compress_module comp_v_83 (
                                            .x(v[83]),
                                            .d(4),
                                            .result(comp_v[83])
                                        );
                                        
                                        compress_module comp_v_84 (
                                            .x(v[84]),
                                            .d(4),
                                            .result(comp_v[84])
                                        );
                                        
                                        compress_module comp_v_85 (
                                            .x(v[85]),
                                            .d(4),
                                            .result(comp_v[85])
                                        );
                                        
                                        compress_module comp_v_86 (
                                            .x(v[86]),
                                            .d(4),
                                            .result(comp_v[86])
                                        );
                                        
                                        compress_module comp_v_87 (
                                            .x(v[87]),
                                            .d(4),
                                            .result(comp_v[87])
                                        );
                                        
                                        compress_module comp_v_88 (
                                            .x(v[88]),
                                            .d(4),
                                            .result(comp_v[88])
                                        );
                                        
                                        compress_module comp_v_89 (
                                            .x(v[89]),
                                            .d(4),
                                            .result(comp_v[89])
                                        );
                                        
                                        compress_module comp_v_90 (
                                            .x(v[90]),
                                            .d(4),
                                            .result(comp_v[90])
                                        );
                                        
                                        compress_module comp_v_91 (
                                            .x(v[91]),
                                            .d(4),
                                            .result(comp_v[91])
                                        );
                                        
                                        compress_module comp_v_92 (
                                            .x(v[92]),
                                            .d(4),
                                            .result(comp_v[92])
                                        );
                                        
                                        compress_module comp_v_93 (
                                            .x(v[93]),
                                            .d(4),
                                            .result(comp_v[93])
                                        );
                                        
                                        compress_module comp_v_94 (
                                            .x(v[94]),
                                            .d(4),
                                            .result(comp_v[94])
                                        );
                                        
                                        compress_module comp_v_95 (
                                            .x(v[95]),
                                            .d(4),
                                            .result(comp_v[95])
                                        );
                                        
                                        compress_module comp_v_96 (
                                            .x(v[96]),
                                            .d(4),
                                            .result(comp_v[96])
                                        );
                                        
                                        compress_module comp_v_97 (
                                            .x(v[97]),
                                            .d(4),
                                            .result(comp_v[97])
                                        );
                                        
                                        compress_module comp_v_98 (
                                            .x(v[98]),
                                            .d(4),
                                            .result(comp_v[98])
                                        );
                                        
                                        compress_module comp_v_99 (
                                            .x(v[99]),
                                            .d(4),
                                            .result(comp_v[99])
                                        );
                                        
                                        compress_module comp_v_100 (
                                            .x(v[100]),
                                            .d(4),
                                            .result(comp_v[100])
                                        );
                                        
                                        compress_module comp_v_101 (
                                            .x(v[101]),
                                            .d(4),
                                            .result(comp_v[101])
                                        );
                                        
                                        compress_module comp_v_102 (
                                            .x(v[102]),
                                            .d(4),
                                            .result(comp_v[102])
                                        );
                                        
                                        compress_module comp_v_103 (
                                            .x(v[103]),
                                            .d(4),
                                            .result(comp_v[103])
                                        );
                                        
                                        compress_module comp_v_104 (
                                            .x(v[104]),
                                            .d(4),
                                            .result(comp_v[104])
                                        );
                                        
                                        compress_module comp_v_105 (
                                            .x(v[105]),
                                            .d(4),
                                            .result(comp_v[105])
                                        );
                                        
                                        compress_module comp_v_106 (
                                            .x(v[106]),
                                            .d(4),
                                            .result(comp_v[106])
                                        );
                                        
                                        compress_module comp_v_107 (
                                            .x(v[107]),
                                            .d(4),
                                            .result(comp_v[107])
                                        );
                                        
                                        compress_module comp_v_108 (
                                            .x(v[108]),
                                            .d(4),
                                            .result(comp_v[108])
                                        );
                                        
                                        compress_module comp_v_109 (
                                            .x(v[109]),
                                            .d(4),
                                            .result(comp_v[109])
                                        );
                                        
                                        compress_module comp_v_110 (
                                            .x(v[110]),
                                            .d(4),
                                            .result(comp_v[110])
                                        );
                                        
                                        compress_module comp_v_111 (
                                            .x(v[111]),
                                            .d(4),
                                            .result(comp_v[111])
                                        );
                                        
                                        compress_module comp_v_112 (
                                            .x(v[112]),
                                            .d(4),
                                            .result(comp_v[112])
                                        );
                                        
                                        compress_module comp_v_113 (
                                            .x(v[113]),
                                            .d(4),
                                            .result(comp_v[113])
                                        );
                                        
                                        compress_module comp_v_114 (
                                            .x(v[114]),
                                            .d(4),
                                            .result(comp_v[114])
                                        );
                                        
                                        compress_module comp_v_115 (
                                            .x(v[115]),
                                            .d(4),
                                            .result(comp_v[115])
                                        );
                                        
                                        compress_module comp_v_116 (
                                            .x(v[116]),
                                            .d(4),
                                            .result(comp_v[116])
                                        );
                                        
                                        compress_module comp_v_117 (
                                            .x(v[117]),
                                            .d(4),
                                            .result(comp_v[117])
                                        );
                                        
                                        compress_module comp_v_118 (
                                            .x(v[118]),
                                            .d(4),
                                            .result(comp_v[118])
                                        );
                                        
                                        compress_module comp_v_119 (
                                            .x(v[119]),
                                            .d(4),
                                            .result(comp_v[119])
                                        );
                                        
                                        compress_module comp_v_120 (
                                            .x(v[120]),
                                            .d(4),
                                            .result(comp_v[120])
                                        );
                                        
                                        compress_module comp_v_121 (
                                            .x(v[121]),
                                            .d(4),
                                            .result(comp_v[121])
                                        );
                                        
                                        compress_module comp_v_122 (
                                            .x(v[122]),
                                            .d(4),
                                            .result(comp_v[122])
                                        );
                                        
                                        compress_module comp_v_123 (
                                            .x(v[123]),
                                            .d(4),
                                            .result(comp_v[123])
                                        );
                                        
                                        compress_module comp_v_124 (
                                            .x(v[124]),
                                            .d(4),
                                            .result(comp_v[124])
                                        );
                                        
                                        compress_module comp_v_125 (
                                            .x(v[125]),
                                            .d(4),
                                            .result(comp_v[125])
                                        );
                                        
                                        compress_module comp_v_126 (
                                            .x(v[126]),
                                            .d(4),
                                            .result(comp_v[126])
                                        );
                                        
                                        compress_module comp_v_127 (
                                            .x(v[127]),
                                            .d(4),
                                            .result(comp_v[127])
                                        );
                                        
                                        compress_module comp_v_128 (
                                            .x(v[128]),
                                            .d(4),
                                            .result(comp_v[128])
                                        );
                                        
                                        compress_module comp_v_129 (
                                            .x(v[129]),
                                            .d(4),
                                            .result(comp_v[129])
                                        );
                                        
                                        compress_module comp_v_130 (
                                            .x(v[130]),
                                            .d(4),
                                            .result(comp_v[130])
                                        );
                                        
                                        compress_module comp_v_131 (
                                            .x(v[131]),
                                            .d(4),
                                            .result(comp_v[131])
                                        );
                                        
                                        compress_module comp_v_132 (
                                            .x(v[132]),
                                            .d(4),
                                            .result(comp_v[132])
                                        );
                                        
                                        compress_module comp_v_133 (
                                            .x(v[133]),
                                            .d(4),
                                            .result(comp_v[133])
                                        );
                                        
                                        compress_module comp_v_134 (
                                            .x(v[134]),
                                            .d(4),
                                            .result(comp_v[134])
                                        );
                                        
                                        compress_module comp_v_135 (
                                            .x(v[135]),
                                            .d(4),
                                            .result(comp_v[135])
                                        );
                                        
                                        compress_module comp_v_136 (
                                            .x(v[136]),
                                            .d(4),
                                            .result(comp_v[136])
                                        );
                                        
                                        compress_module comp_v_137 (
                                            .x(v[137]),
                                            .d(4),
                                            .result(comp_v[137])
                                        );
                                        
                                        compress_module comp_v_138 (
                                            .x(v[138]),
                                            .d(4),
                                            .result(comp_v[138])
                                        );
                                        
                                        compress_module comp_v_139 (
                                            .x(v[139]),
                                            .d(4),
                                            .result(comp_v[139])
                                        );
                                        
                                        compress_module comp_v_140 (
                                            .x(v[140]),
                                            .d(4),
                                            .result(comp_v[140])
                                        );
                                        
                                        compress_module comp_v_141 (
                                            .x(v[141]),
                                            .d(4),
                                            .result(comp_v[141])
                                        );
                                        
                                        compress_module comp_v_142 (
                                            .x(v[142]),
                                            .d(4),
                                            .result(comp_v[142])
                                        );
                                        
                                        compress_module comp_v_143 (
                                            .x(v[143]),
                                            .d(4),
                                            .result(comp_v[143])
                                        );
                                        
                                        compress_module comp_v_144 (
                                            .x(v[144]),
                                            .d(4),
                                            .result(comp_v[144])
                                        );
                                        
                                        compress_module comp_v_145 (
                                            .x(v[145]),
                                            .d(4),
                                            .result(comp_v[145])
                                        );
                                        
                                        compress_module comp_v_146 (
                                            .x(v[146]),
                                            .d(4),
                                            .result(comp_v[146])
                                        );
                                        
                                        compress_module comp_v_147 (
                                            .x(v[147]),
                                            .d(4),
                                            .result(comp_v[147])
                                        );
                                        
                                        compress_module comp_v_148 (
                                            .x(v[148]),
                                            .d(4),
                                            .result(comp_v[148])
                                        );
                                        
                                        compress_module comp_v_149 (
                                            .x(v[149]),
                                            .d(4),
                                            .result(comp_v[149])
                                        );
                                        
                                        compress_module comp_v_150 (
                                            .x(v[150]),
                                            .d(4),
                                            .result(comp_v[150])
                                        );
                                        
                                        compress_module comp_v_151 (
                                            .x(v[151]),
                                            .d(4),
                                            .result(comp_v[151])
                                        );
                                        
                                        compress_module comp_v_152 (
                                            .x(v[152]),
                                            .d(4),
                                            .result(comp_v[152])
                                        );
                                        
                                        compress_module comp_v_153 (
                                            .x(v[153]),
                                            .d(4),
                                            .result(comp_v[153])
                                        );
                                        
                                        compress_module comp_v_154 (
                                            .x(v[154]),
                                            .d(4),
                                            .result(comp_v[154])
                                        );
                                        
                                        compress_module comp_v_155 (
                                            .x(v[155]),
                                            .d(4),
                                            .result(comp_v[155])
                                        );
                                        
                                        compress_module comp_v_156 (
                                            .x(v[156]),
                                            .d(4),
                                            .result(comp_v[156])
                                        );
                                        
                                        compress_module comp_v_157 (
                                            .x(v[157]),
                                            .d(4),
                                            .result(comp_v[157])
                                        );
                                        
                                        compress_module comp_v_158 (
                                            .x(v[158]),
                                            .d(4),
                                            .result(comp_v[158])
                                        );
                                        
                                        compress_module comp_v_159 (
                                            .x(v[159]),
                                            .d(4),
                                            .result(comp_v[159])
                                        );
                                        
                                        compress_module comp_v_160 (
                                            .x(v[160]),
                                            .d(4),
                                            .result(comp_v[160])
                                        );
                                        
                                        compress_module comp_v_161 (
                                            .x(v[161]),
                                            .d(4),
                                            .result(comp_v[161])
                                        );
                                        
                                        compress_module comp_v_162 (
                                            .x(v[162]),
                                            .d(4),
                                            .result(comp_v[162])
                                        );
                                        
                                        compress_module comp_v_163 (
                                            .x(v[163]),
                                            .d(4),
                                            .result(comp_v[163])
                                        );
                                        
                                        compress_module comp_v_164 (
                                            .x(v[164]),
                                            .d(4),
                                            .result(comp_v[164])
                                        );
                                        
                                        compress_module comp_v_165 (
                                            .x(v[165]),
                                            .d(4),
                                            .result(comp_v[165])
                                        );
                                        
                                        compress_module comp_v_166 (
                                            .x(v[166]),
                                            .d(4),
                                            .result(comp_v[166])
                                        );
                                        
                                        compress_module comp_v_167 (
                                            .x(v[167]),
                                            .d(4),
                                            .result(comp_v[167])
                                        );
                                        
                                        compress_module comp_v_168 (
                                            .x(v[168]),
                                            .d(4),
                                            .result(comp_v[168])
                                        );
                                        
                                        compress_module comp_v_169 (
                                            .x(v[169]),
                                            .d(4),
                                            .result(comp_v[169])
                                        );
                                        
                                        compress_module comp_v_170 (
                                            .x(v[170]),
                                            .d(4),
                                            .result(comp_v[170])
                                        );
                                        
                                        compress_module comp_v_171 (
                                            .x(v[171]),
                                            .d(4),
                                            .result(comp_v[171])
                                        );
                                        
                                        compress_module comp_v_172 (
                                            .x(v[172]),
                                            .d(4),
                                            .result(comp_v[172])
                                        );
                                        
                                        compress_module comp_v_173 (
                                            .x(v[173]),
                                            .d(4),
                                            .result(comp_v[173])
                                        );
                                        
                                        compress_module comp_v_174 (
                                            .x(v[174]),
                                            .d(4),
                                            .result(comp_v[174])
                                        );
                                        
                                        compress_module comp_v_175 (
                                            .x(v[175]),
                                            .d(4),
                                            .result(comp_v[175])
                                        );
                                        
                                        compress_module comp_v_176 (
                                            .x(v[176]),
                                            .d(4),
                                            .result(comp_v[176])
                                        );
                                        
                                        compress_module comp_v_177 (
                                            .x(v[177]),
                                            .d(4),
                                            .result(comp_v[177])
                                        );
                                        
                                        compress_module comp_v_178 (
                                            .x(v[178]),
                                            .d(4),
                                            .result(comp_v[178])
                                        );
                                        
                                        compress_module comp_v_179 (
                                            .x(v[179]),
                                            .d(4),
                                            .result(comp_v[179])
                                        );
                                        
                                        compress_module comp_v_180 (
                                            .x(v[180]),
                                            .d(4),
                                            .result(comp_v[180])
                                        );
                                        
                                        compress_module comp_v_181 (
                                            .x(v[181]),
                                            .d(4),
                                            .result(comp_v[181])
                                        );
                                        
                                        compress_module comp_v_182 (
                                            .x(v[182]),
                                            .d(4),
                                            .result(comp_v[182])
                                        );
                                        
                                        compress_module comp_v_183 (
                                            .x(v[183]),
                                            .d(4),
                                            .result(comp_v[183])
                                        );
                                        
                                        compress_module comp_v_184 (
                                            .x(v[184]),
                                            .d(4),
                                            .result(comp_v[184])
                                        );
                                        
                                        compress_module comp_v_185 (
                                            .x(v[185]),
                                            .d(4),
                                            .result(comp_v[185])
                                        );
                                        
                                        compress_module comp_v_186 (
                                            .x(v[186]),
                                            .d(4),
                                            .result(comp_v[186])
                                        );
                                        
                                        compress_module comp_v_187 (
                                            .x(v[187]),
                                            .d(4),
                                            .result(comp_v[187])
                                        );
                                        
                                        compress_module comp_v_188 (
                                            .x(v[188]),
                                            .d(4),
                                            .result(comp_v[188])
                                        );
                                        
                                        compress_module comp_v_189 (
                                            .x(v[189]),
                                            .d(4),
                                            .result(comp_v[189])
                                        );
                                        
                                        compress_module comp_v_190 (
                                            .x(v[190]),
                                            .d(4),
                                            .result(comp_v[190])
                                        );
                                        
                                        compress_module comp_v_191 (
                                            .x(v[191]),
                                            .d(4),
                                            .result(comp_v[191])
                                        );
                                        
                                        compress_module comp_v_192 (
                                            .x(v[192]),
                                            .d(4),
                                            .result(comp_v[192])
                                        );
                                        
                                        compress_module comp_v_193 (
                                            .x(v[193]),
                                            .d(4),
                                            .result(comp_v[193])
                                        );
                                        
                                        compress_module comp_v_194 (
                                            .x(v[194]),
                                            .d(4),
                                            .result(comp_v[194])
                                        );
                                        
                                        compress_module comp_v_195 (
                                            .x(v[195]),
                                            .d(4),
                                            .result(comp_v[195])
                                        );
                                        
                                        compress_module comp_v_196 (
                                            .x(v[196]),
                                            .d(4),
                                            .result(comp_v[196])
                                        );
                                        
                                        compress_module comp_v_197 (
                                            .x(v[197]),
                                            .d(4),
                                            .result(comp_v[197])
                                        );
                                        
                                        compress_module comp_v_198 (
                                            .x(v[198]),
                                            .d(4),
                                            .result(comp_v[198])
                                        );
                                        
                                        compress_module comp_v_199 (
                                            .x(v[199]),
                                            .d(4),
                                            .result(comp_v[199])
                                        );
                                        
                                        compress_module comp_v_200 (
                                            .x(v[200]),
                                            .d(4),
                                            .result(comp_v[200])
                                        );
                                        
                                        compress_module comp_v_201 (
                                            .x(v[201]),
                                            .d(4),
                                            .result(comp_v[201])
                                        );
                                        
                                        compress_module comp_v_202 (
                                            .x(v[202]),
                                            .d(4),
                                            .result(comp_v[202])
                                        );
                                        
                                        compress_module comp_v_203 (
                                            .x(v[203]),
                                            .d(4),
                                            .result(comp_v[203])
                                        );
                                        
                                        compress_module comp_v_204 (
                                            .x(v[204]),
                                            .d(4),
                                            .result(comp_v[204])
                                        );
                                        
                                        compress_module comp_v_205 (
                                            .x(v[205]),
                                            .d(4),
                                            .result(comp_v[205])
                                        );
                                        
                                        compress_module comp_v_206 (
                                            .x(v[206]),
                                            .d(4),
                                            .result(comp_v[206])
                                        );
                                        
                                        compress_module comp_v_207 (
                                            .x(v[207]),
                                            .d(4),
                                            .result(comp_v[207])
                                        );
                                        
                                        compress_module comp_v_208 (
                                            .x(v[208]),
                                            .d(4),
                                            .result(comp_v[208])
                                        );
                                        
                                        compress_module comp_v_209 (
                                            .x(v[209]),
                                            .d(4),
                                            .result(comp_v[209])
                                        );
                                        
                                        compress_module comp_v_210 (
                                            .x(v[210]),
                                            .d(4),
                                            .result(comp_v[210])
                                        );
                                        
                                        compress_module comp_v_211 (
                                            .x(v[211]),
                                            .d(4),
                                            .result(comp_v[211])
                                        );
                                        
                                        compress_module comp_v_212 (
                                            .x(v[212]),
                                            .d(4),
                                            .result(comp_v[212])
                                        );
                                        
                                        compress_module comp_v_213 (
                                            .x(v[213]),
                                            .d(4),
                                            .result(comp_v[213])
                                        );
                                        
                                        compress_module comp_v_214 (
                                            .x(v[214]),
                                            .d(4),
                                            .result(comp_v[214])
                                        );
                                        
                                        compress_module comp_v_215 (
                                            .x(v[215]),
                                            .d(4),
                                            .result(comp_v[215])
                                        );
                                        
                                        compress_module comp_v_216 (
                                            .x(v[216]),
                                            .d(4),
                                            .result(comp_v[216])
                                        );
                                        
                                        compress_module comp_v_217 (
                                            .x(v[217]),
                                            .d(4),
                                            .result(comp_v[217])
                                        );
                                        
                                        compress_module comp_v_218 (
                                            .x(v[218]),
                                            .d(4),
                                            .result(comp_v[218])
                                        );
                                        
                                        compress_module comp_v_219 (
                                            .x(v[219]),
                                            .d(4),
                                            .result(comp_v[219])
                                        );
                                        
                                        compress_module comp_v_220 (
                                            .x(v[220]),
                                            .d(4),
                                            .result(comp_v[220])
                                        );
                                        
                                        compress_module comp_v_221 (
                                            .x(v[221]),
                                            .d(4),
                                            .result(comp_v[221])
                                        );
                                        
                                        compress_module comp_v_222 (
                                            .x(v[222]),
                                            .d(4),
                                            .result(comp_v[222])
                                        );
                                        
                                        compress_module comp_v_223 (
                                            .x(v[223]),
                                            .d(4),
                                            .result(comp_v[223])
                                        );
                                        
                                        compress_module comp_v_224 (
                                            .x(v[224]),
                                            .d(4),
                                            .result(comp_v[224])
                                        );
                                        
                                        compress_module comp_v_225 (
                                            .x(v[225]),
                                            .d(4),
                                            .result(comp_v[225])
                                        );
                                        
                                        compress_module comp_v_226 (
                                            .x(v[226]),
                                            .d(4),
                                            .result(comp_v[226])
                                        );
                                        
                                        compress_module comp_v_227 (
                                            .x(v[227]),
                                            .d(4),
                                            .result(comp_v[227])
                                        );
                                        
                                        compress_module comp_v_228 (
                                            .x(v[228]),
                                            .d(4),
                                            .result(comp_v[228])
                                        );
                                        
                                        compress_module comp_v_229 (
                                            .x(v[229]),
                                            .d(4),
                                            .result(comp_v[229])
                                        );
                                        
                                        compress_module comp_v_230 (
                                            .x(v[230]),
                                            .d(4),
                                            .result(comp_v[230])
                                        );
                                        
                                        compress_module comp_v_231 (
                                            .x(v[231]),
                                            .d(4),
                                            .result(comp_v[231])
                                        );
                                        
                                        compress_module comp_v_232 (
                                            .x(v[232]),
                                            .d(4),
                                            .result(comp_v[232])
                                        );
                                        
                                        compress_module comp_v_233 (
                                            .x(v[233]),
                                            .d(4),
                                            .result(comp_v[233])
                                        );
                                        
                                        compress_module comp_v_234 (
                                            .x(v[234]),
                                            .d(4),
                                            .result(comp_v[234])
                                        );
                                        
                                        compress_module comp_v_235 (
                                            .x(v[235]),
                                            .d(4),
                                            .result(comp_v[235])
                                        );
                                        
                                        compress_module comp_v_236 (
                                            .x(v[236]),
                                            .d(4),
                                            .result(comp_v[236])
                                        );
                                        
                                        compress_module comp_v_237 (
                                            .x(v[237]),
                                            .d(4),
                                            .result(comp_v[237])
                                        );
                                        
                                        compress_module comp_v_238 (
                                            .x(v[238]),
                                            .d(4),
                                            .result(comp_v[238])
                                        );
                                        
                                        compress_module comp_v_239 (
                                            .x(v[239]),
                                            .d(4),
                                            .result(comp_v[239])
                                        );
                                        
                                        compress_module comp_v_240 (
                                            .x(v[240]),
                                            .d(4),
                                            .result(comp_v[240])
                                        );
                                        
                                        compress_module comp_v_241 (
                                            .x(v[241]),
                                            .d(4),
                                            .result(comp_v[241])
                                        );
                                        
                                        compress_module comp_v_242 (
                                            .x(v[242]),
                                            .d(4),
                                            .result(comp_v[242])
                                        );
                                        
                                        compress_module comp_v_243 (
                                            .x(v[243]),
                                            .d(4),
                                            .result(comp_v[243])
                                        );
                                        
                                        compress_module comp_v_244 (
                                            .x(v[244]),
                                            .d(4),
                                            .result(comp_v[244])
                                        );
                                        
                                        compress_module comp_v_245 (
                                            .x(v[245]),
                                            .d(4),
                                            .result(comp_v[245])
                                        );
                                        
                                        compress_module comp_v_246 (
                                            .x(v[246]),
                                            .d(4),
                                            .result(comp_v[246])
                                        );
                                        
                                        compress_module comp_v_247 (
                                            .x(v[247]),
                                            .d(4),
                                            .result(comp_v[247])
                                        );
                                        
                                        compress_module comp_v_248 (
                                            .x(v[248]),
                                            .d(4),
                                            .result(comp_v[248])
                                        );
                                        
                                        compress_module comp_v_249 (
                                            .x(v[249]),
                                            .d(4),
                                            .result(comp_v[249])
                                        );
                                        
                                        compress_module comp_v_250 (
                                            .x(v[250]),
                                            .d(4),
                                            .result(comp_v[250])
                                        );
                                        
                                        compress_module comp_v_251 (
                                            .x(v[251]),
                                            .d(4),
                                            .result(comp_v[251])
                                        );
                                        
                                        compress_module comp_v_252 (
                                            .x(v[252]),
                                            .d(4),
                                            .result(comp_v[252])
                                        );
                                        
                                        compress_module comp_v_253 (
                                            .x(v[253]),
                                            .d(4),
                                            .result(comp_v[253])
                                        );
                                        
                                        compress_module comp_v_254 (
                                            .x(v[254]),
                                            .d(4),
                                            .result(comp_v[254])
                                        );
                                        
                                        compress_module comp_v_255 (
                                            .x(v[255]),
                                            .d(4),
                                            .result(comp_v[255])
                                        );
                                        encode #(.D(8),.BYTE_LEN(32))enc_u0 (
                                            .F(com_out[0]),
                                            .B(encode_u[0])
                                        );
                                        
                                        encode #(.D(8),.BYTE_LEN(32))enc_u1 (
                                            .F(com_out[1]),
                                            .B(encode_u[1])
                                        );
                                        
                                        encode #(.D(8),.BYTE_LEN(32))enc_u2 (
                                            .F(com_out[2]),
                                            .B(encode_u[2])
                                        );
                                       encode #(.D(4),.BYTE_LEN(32))enc_v0 (
                                            .F(comp_v[0]),
                                            .B(encode_v[0])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v1 (
                                            .F(comp_v[1]),
                                            .B(encode_v[1])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v2 (
                                            .F(comp_v[2]),
                                            .B(encode_v[2])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v3 (
                                            .F(comp_v[3]),
                                            .B(encode_v[3])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v4 (
                                            .F(comp_v[4]),
                                            .B(encode_v[4])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v5 (
                                            .F(comp_v[5]),
                                            .B(encode_v[5])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v6 (
                                            .F(comp_v[6]),
                                            .B(encode_v[6])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v7 (
                                            .F(comp_v[7]),
                                            .B(encode_v[7])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v8 (
                                            .F(comp_v[8]),
                                            .B(encode_v[8])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v9 (
                                            .F(comp_v[9]),
                                            .B(encode_v[9])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v10 (
                                            .F(comp_v[10]),
                                            .B(encode_v[10])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v11 (
                                            .F(comp_v[11]),
                                            .B(encode_v[11])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v12 (
                                            .F(comp_v[12]),
                                            .B(encode_v[12])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v13 (
                                            .F(comp_v[13]),
                                            .B(encode_v[13])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v14 (
                                            .F(comp_v[14]),
                                            .B(encode_v[14])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v15 (
                                            .F(comp_v[15]),
                                            .B(encode_v[15])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v16 (
                                            .F(comp_v[16]),
                                            .B(encode_v[16])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v17 (
                                            .F(comp_v[17]),
                                            .B(encode_v[17])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v18 (
                                            .F(comp_v[18]),
                                            .B(encode_v[18])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v19 (
                                            .F(comp_v[19]),
                                            .B(encode_v[19])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v20 (
                                            .F(comp_v[20]),
                                            .B(encode_v[20])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v21 (
                                            .F(comp_v[21]),
                                            .B(encode_v[21])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v22 (
                                            .F(comp_v[22]),
                                            .B(encode_v[22])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v23 (
                                            .F(comp_v[23]),
                                            .B(encode_v[23])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v24 (
                                            .F(comp_v[24]),
                                            .B(encode_v[24])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v25 (
                                            .F(comp_v[25]),
                                            .B(encode_v[25])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v26 (
                                            .F(comp_v[26]),
                                            .B(encode_v[26])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v27 (
                                            .F(comp_v[27]),
                                            .B(encode_v[27])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v28 (
                                            .F(comp_v[28]),
                                            .B(encode_v[28])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v29 (
                                            .F(comp_v[29]),
                                            .B(encode_v[29])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v30 (
                                            .F(comp_v[30]),
                                            .B(encode_v[30])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v31 (
                                            .F(comp_v[31]),
                                            .B(encode_v[31])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v32 (
                                            .F(comp_v[32]),
                                            .B(encode_v[32])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v33 (
                                            .F(comp_v[33]),
                                            .B(encode_v[33])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v34 (
                                            .F(comp_v[34]),
                                            .B(encode_v[34])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v35 (
                                            .F(comp_v[35]),
                                            .B(encode_v[35])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v36 (
                                            .F(comp_v[36]),
                                            .B(encode_v[36])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v37 (
                                            .F(comp_v[37]),
                                            .B(encode_v[37])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v38 (
                                            .F(comp_v[38]),
                                            .B(encode_v[38])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v39 (
                                            .F(comp_v[39]),
                                            .B(encode_v[39])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v40 (
                                            .F(comp_v[40]),
                                            .B(encode_v[40])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v41 (
                                            .F(comp_v[41]),
                                            .B(encode_v[41])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v42 (
                                            .F(comp_v[42]),
                                            .B(encode_v[42])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v43 (
                                            .F(comp_v[43]),
                                            .B(encode_v[43])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v44 (
                                            .F(comp_v[44]),
                                            .B(encode_v[44])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v45 (
                                            .F(comp_v[45]),
                                            .B(encode_v[45])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v46 (
                                            .F(comp_v[46]),
                                            .B(encode_v[46])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v47 (
                                            .F(comp_v[47]),
                                            .B(encode_v[47])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v48 (
                                            .F(comp_v[48]),
                                            .B(encode_v[48])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v49 (
                                            .F(comp_v[49]),
                                            .B(encode_v[49])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v50 (
                                            .F(comp_v[50]),
                                            .B(encode_v[50])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v51 (
                                            .F(comp_v[51]),
                                            .B(encode_v[51])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v52 (
                                            .F(comp_v[52]),
                                            .B(encode_v[52])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v53 (
                                            .F(comp_v[53]),
                                            .B(encode_v[53])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v54 (
                                            .F(comp_v[54]),
                                            .B(encode_v[54])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v55 (
                                            .F(comp_v[55]),
                                            .B(encode_v[55])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v56 (
                                            .F(comp_v[56]),
                                            .B(encode_v[56])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v57 (
                                            .F(comp_v[57]),
                                            .B(encode_v[57])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v58 (
                                            .F(comp_v[58]),
                                            .B(encode_v[58])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v59 (
                                            .F(comp_v[59]),
                                            .B(encode_v[59])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v60 (
                                            .F(comp_v[60]),
                                            .B(encode_v[60])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v61 (
                                            .F(comp_v[61]),
                                            .B(encode_v[61])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v62 (
                                            .F(comp_v[62]),
                                            .B(encode_v[62])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v63 (
                                            .F(comp_v[63]),
                                            .B(encode_v[63])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v64 (
                                            .F(comp_v[64]),
                                            .B(encode_v[64])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v65 (
                                            .F(comp_v[65]),
                                            .B(encode_v[65])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v66 (
                                            .F(comp_v[66]),
                                            .B(encode_v[66])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v67 (
                                            .F(comp_v[67]),
                                            .B(encode_v[67])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v68 (
                                            .F(comp_v[68]),
                                            .B(encode_v[68])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v69 (
                                            .F(comp_v[69]),
                                            .B(encode_v[69])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v70 (
                                            .F(comp_v[70]),
                                            .B(encode_v[70])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v71 (
                                            .F(comp_v[71]),
                                            .B(encode_v[71])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v72 (
                                            .F(comp_v[72]),
                                            .B(encode_v[72])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v73 (
                                            .F(comp_v[73]),
                                            .B(encode_v[73])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v74 (
                                            .F(comp_v[74]),
                                            .B(encode_v[74])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v75 (
                                            .F(comp_v[75]),
                                            .B(encode_v[75])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v76 (
                                            .F(comp_v[76]),
                                            .B(encode_v[76])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v77 (
                                            .F(comp_v[77]),
                                            .B(encode_v[77])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v78 (
                                            .F(comp_v[78]),
                                            .B(encode_v[78])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v79 (
                                            .F(comp_v[79]),
                                            .B(encode_v[79])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v80 (
                                            .F(comp_v[80]),
                                            .B(encode_v[80])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v81 (
                                            .F(comp_v[81]),
                                            .B(encode_v[81])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v82 (
                                            .F(comp_v[82]),
                                            .B(encode_v[82])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v83 (
                                            .F(comp_v[83]),
                                            .B(encode_v[83])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v84 (
                                            .F(comp_v[84]),
                                            .B(encode_v[84])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v85 (
                                            .F(comp_v[85]),
                                            .B(encode_v[85])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v86 (
                                            .F(comp_v[86]),
                                            .B(encode_v[86])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v87 (
                                            .F(comp_v[87]),
                                            .B(encode_v[87])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v88 (
                                            .F(comp_v[88]),
                                            .B(encode_v[88])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v89 (
                                            .F(comp_v[89]),
                                            .B(encode_v[89])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v90 (
                                            .F(comp_v[90]),
                                            .B(encode_v[90])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v91 (
                                            .F(comp_v[91]),
                                            .B(encode_v[91])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v92 (
                                            .F(comp_v[92]),
                                            .B(encode_v[92])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v93 (
                                            .F(comp_v[93]),
                                            .B(encode_v[93])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v94 (
                                            .F(comp_v[94]),
                                            .B(encode_v[94])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v95 (
                                            .F(comp_v[95]),
                                            .B(encode_v[95])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v96 (
                                            .F(comp_v[96]),
                                            .B(encode_v[96])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v97 (
                                            .F(comp_v[97]),
                                            .B(encode_v[97])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v98 (
                                            .F(comp_v[98]),
                                            .B(encode_v[98])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v99 (
                                            .F(comp_v[99]),
                                            .B(encode_v[99])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v100 (
                                            .F(comp_v[100]),
                                            .B(encode_v[100])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v101 (
                                            .F(comp_v[101]),
                                            .B(encode_v[101])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v102 (
                                            .F(comp_v[102]),
                                            .B(encode_v[102])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v103 (
                                            .F(comp_v[103]),
                                            .B(encode_v[103])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v104 (
                                            .F(comp_v[104]),
                                            .B(encode_v[104])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v105 (
                                            .F(comp_v[105]),
                                            .B(encode_v[105])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v106 (
                                            .F(comp_v[106]),
                                            .B(encode_v[106])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v107 (
                                            .F(comp_v[107]),
                                            .B(encode_v[107])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v108 (
                                            .F(comp_v[108]),
                                            .B(encode_v[108])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v109 (
                                            .F(comp_v[109]),
                                            .B(encode_v[109])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v110 (
                                            .F(comp_v[110]),
                                            .B(encode_v[110])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v111 (
                                            .F(comp_v[111]),
                                            .B(encode_v[111])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v112 (
                                            .F(comp_v[112]),
                                            .B(encode_v[112])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v113 (
                                            .F(comp_v[113]),
                                            .B(encode_v[113])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v114 (
                                            .F(comp_v[114]),
                                            .B(encode_v[114])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v115 (
                                            .F(comp_v[115]),
                                            .B(encode_v[115])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v116 (
                                            .F(comp_v[116]),
                                            .B(encode_v[116])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v117 (
                                            .F(comp_v[117]),
                                            .B(encode_v[117])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v118 (
                                            .F(comp_v[118]),
                                            .B(encode_v[118])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v119 (
                                            .F(comp_v[119]),
                                            .B(encode_v[119])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v120 (
                                            .F(comp_v[120]),
                                            .B(encode_v[120])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v121 (
                                            .F(comp_v[121]),
                                            .B(encode_v[121])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v122 (
                                            .F(comp_v[122]),
                                            .B(encode_v[122])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v123 (
                                            .F(comp_v[123]),
                                            .B(encode_v[123])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v124 (
                                            .F(comp_v[124]),
                                            .B(encode_v[124])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v125 (
                                            .F(comp_v[125]),
                                            .B(encode_v[125])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v126 (
                                            .F(comp_v[126]),
                                            .B(encode_v[126])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v127 (
                                            .F(comp_v[127]),
                                            .B(encode_v[127])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v128 (
                                            .F(comp_v[128]),
                                            .B(encode_v[128])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v129 (
                                            .F(comp_v[129]),
                                            .B(encode_v[129])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v130 (
                                            .F(comp_v[130]),
                                            .B(encode_v[130])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v131 (
                                            .F(comp_v[131]),
                                            .B(encode_v[131])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v132 (
                                            .F(comp_v[132]),
                                            .B(encode_v[132])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v133 (
                                            .F(comp_v[133]),
                                            .B(encode_v[133])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v134 (
                                            .F(comp_v[134]),
                                            .B(encode_v[134])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v135 (
                                            .F(comp_v[135]),
                                            .B(encode_v[135])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v136 (
                                            .F(comp_v[136]),
                                            .B(encode_v[136])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v137 (
                                            .F(comp_v[137]),
                                            .B(encode_v[137])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v138 (
                                            .F(comp_v[138]),
                                            .B(encode_v[138])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v139 (
                                            .F(comp_v[139]),
                                            .B(encode_v[139])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v140 (
                                            .F(comp_v[140]),
                                            .B(encode_v[140])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v141 (
                                            .F(comp_v[141]),
                                            .B(encode_v[141])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v142 (
                                            .F(comp_v[142]),
                                            .B(encode_v[142])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v143 (
                                            .F(comp_v[143]),
                                            .B(encode_v[143])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v144 (
                                            .F(comp_v[144]),
                                            .B(encode_v[144])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v145 (
                                            .F(comp_v[145]),
                                            .B(encode_v[145])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v146 (
                                            .F(comp_v[146]),
                                            .B(encode_v[146])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v147 (
                                            .F(comp_v[147]),
                                            .B(encode_v[147])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v148 (
                                            .F(comp_v[148]),
                                            .B(encode_v[148])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v149 (
                                            .F(comp_v[149]),
                                            .B(encode_v[149])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v150 (
                                            .F(comp_v[150]),
                                            .B(encode_v[150])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v151 (
                                            .F(comp_v[151]),
                                            .B(encode_v[151])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v152 (
                                            .F(comp_v[152]),
                                            .B(encode_v[152])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v153 (
                                            .F(comp_v[153]),
                                            .B(encode_v[153])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v154 (
                                            .F(comp_v[154]),
                                            .B(encode_v[154])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v155 (
                                            .F(comp_v[155]),
                                            .B(encode_v[155])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v156 (
                                            .F(comp_v[156]),
                                            .B(encode_v[156])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v157 (
                                            .F(comp_v[157]),
                                            .B(encode_v[157])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v158 (
                                            .F(comp_v[158]),
                                            .B(encode_v[158])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v159 (
                                            .F(comp_v[159]),
                                            .B(encode_v[159])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v160 (
                                            .F(comp_v[160]),
                                            .B(encode_v[160])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v161 (
                                            .F(comp_v[161]),
                                            .B(encode_v[161])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v162 (
                                            .F(comp_v[162]),
                                            .B(encode_v[162])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v163 (
                                            .F(comp_v[163]),
                                            .B(encode_v[163])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v164 (
                                            .F(comp_v[164]),
                                            .B(encode_v[164])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v165 (
                                            .F(comp_v[165]),
                                            .B(encode_v[165])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v166 (
                                            .F(comp_v[166]),
                                            .B(encode_v[166])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v167 (
                                            .F(comp_v[167]),
                                            .B(encode_v[167])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v168 (
                                            .F(comp_v[168]),
                                            .B(encode_v[168])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v169 (
                                            .F(comp_v[169]),
                                            .B(encode_v[169])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v170 (
                                            .F(comp_v[170]),
                                            .B(encode_v[170])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v171 (
                                            .F(comp_v[171]),
                                            .B(encode_v[171])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v172 (
                                            .F(comp_v[172]),
                                            .B(encode_v[172])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v173 (
                                            .F(comp_v[173]),
                                            .B(encode_v[173])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v174 (
                                            .F(comp_v[174]),
                                            .B(encode_v[174])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v175 (
                                            .F(comp_v[175]),
                                            .B(encode_v[175])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v176 (
                                            .F(comp_v[176]),
                                            .B(encode_v[176])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v177 (
                                            .F(comp_v[177]),
                                            .B(encode_v[177])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v178 (
                                            .F(comp_v[178]),
                                            .B(encode_v[178])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v179 (
                                            .F(comp_v[179]),
                                            .B(encode_v[179])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v180 (
                                            .F(comp_v[180]),
                                            .B(encode_v[180])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v181 (
                                            .F(comp_v[181]),
                                            .B(encode_v[181])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v182 (
                                            .F(comp_v[182]),
                                            .B(encode_v[182])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v183 (
                                            .F(comp_v[183]),
                                            .B(encode_v[183])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v184 (
                                            .F(comp_v[184]),
                                            .B(encode_v[184])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v185 (
                                            .F(comp_v[185]),
                                            .B(encode_v[185])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v186 (
                                            .F(comp_v[186]),
                                            .B(encode_v[186])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v187 (
                                            .F(comp_v[187]),
                                            .B(encode_v[187])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v188 (
                                            .F(comp_v[188]),
                                            .B(encode_v[188])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v189 (
                                            .F(comp_v[189]),
                                            .B(encode_v[189])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v190 (
                                            .F(comp_v[190]),
                                            .B(encode_v[190])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v191 (
                                            .F(comp_v[191]),
                                            .B(encode_v[191])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v192 (
                                            .F(comp_v[192]),
                                            .B(encode_v[192])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v193 (
                                            .F(comp_v[193]),
                                            .B(encode_v[193])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v194 (
                                            .F(comp_v[194]),
                                            .B(encode_v[194])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v195 (
                                            .F(comp_v[195]),
                                            .B(encode_v[195])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v196 (
                                            .F(comp_v[196]),
                                            .B(encode_v[196])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v197 (
                                            .F(comp_v[197]),
                                            .B(encode_v[197])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v198 (
                                            .F(comp_v[198]),
                                            .B(encode_v[198])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v199 (
                                            .F(comp_v[199]),
                                            .B(encode_v[199])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v200 (
                                            .F(comp_v[200]),
                                            .B(encode_v[200])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v201 (
                                            .F(comp_v[201]),
                                            .B(encode_v[201])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v202 (
                                            .F(comp_v[202]),
                                            .B(encode_v[202])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v203 (
                                            .F(comp_v[203]),
                                            .B(encode_v[203])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v204 (
                                            .F(comp_v[204]),
                                            .B(encode_v[204])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v205 (
                                            .F(comp_v[205]),
                                            .B(encode_v[205])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v206 (
                                            .F(comp_v[206]),
                                            .B(encode_v[206])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v207 (
                                            .F(comp_v[207]),
                                            .B(encode_v[207])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v208 (
                                            .F(comp_v[208]),
                                            .B(encode_v[208])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v209 (
                                            .F(comp_v[209]),
                                            .B(encode_v[209])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v210 (
                                            .F(comp_v[210]),
                                            .B(encode_v[210])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v211 (
                                            .F(comp_v[211]),
                                            .B(encode_v[211])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v212 (
                                            .F(comp_v[212]),
                                            .B(encode_v[212])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v213 (
                                            .F(comp_v[213]),
                                            .B(encode_v[213])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v214 (
                                            .F(comp_v[214]),
                                            .B(encode_v[214])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v215 (
                                            .F(comp_v[215]),
                                            .B(encode_v[215])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v216 (
                                            .F(comp_v[216]),
                                            .B(encode_v[216])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v217 (
                                            .F(comp_v[217]),
                                            .B(encode_v[217])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v218 (
                                            .F(comp_v[218]),
                                            .B(encode_v[218])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v219 (
                                            .F(comp_v[219]),
                                            .B(encode_v[219])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v220 (
                                            .F(comp_v[220]),
                                            .B(encode_v[220])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v221 (
                                            .F(comp_v[221]),
                                            .B(encode_v[221])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v222 (
                                            .F(comp_v[222]),
                                            .B(encode_v[222])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v223 (
                                            .F(comp_v[223]),
                                            .B(encode_v[223])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v224 (
                                            .F(comp_v[224]),
                                            .B(encode_v[224])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v225 (
                                            .F(comp_v[225]),
                                            .B(encode_v[225])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v226 (
                                            .F(comp_v[226]),
                                            .B(encode_v[226])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v227 (
                                            .F(comp_v[227]),
                                            .B(encode_v[227])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v228 (
                                            .F(comp_v[228]),
                                            .B(encode_v[228])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v229 (
                                            .F(comp_v[229]),
                                            .B(encode_v[229])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v230 (
                                            .F(comp_v[230]),
                                            .B(encode_v[230])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v231 (
                                            .F(comp_v[231]),
                                            .B(encode_v[231])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v232 (
                                            .F(comp_v[232]),
                                            .B(encode_v[232])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v233 (
                                            .F(comp_v[233]),
                                            .B(encode_v[233])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v234 (
                                            .F(comp_v[234]),
                                            .B(encode_v[234])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v235 (
                                            .F(comp_v[235]),
                                            .B(encode_v[235])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v236 (
                                            .F(comp_v[236]),
                                            .B(encode_v[236])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v237 (
                                            .F(comp_v[237]),
                                            .B(encode_v[237])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v238 (
                                            .F(comp_v[238]),
                                            .B(encode_v[238])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v239 (
                                            .F(comp_v[239]),
                                            .B(encode_v[239])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v240 (
                                            .F(comp_v[240]),
                                            .B(encode_v[240])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v241 (
                                            .F(comp_v[241]),
                                            .B(encode_v[241])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v242 (
                                            .F(comp_v[242]),
                                            .B(encode_v[242])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v243 (
                                            .F(comp_v[243]),
                                            .B(encode_v[243])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v244 (
                                            .F(comp_v[244]),
                                            .B(encode_v[244])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v245 (
                                            .F(comp_v[245]),
                                            .B(encode_v[245])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v246 (
                                            .F(comp_v[246]),
                                            .B(encode_v[246])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v247 (
                                            .F(comp_v[247]),
                                            .B(encode_v[247])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v248 (
                                            .F(comp_v[248]),
                                            .B(encode_v[248])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v249 (
                                            .F(comp_v[249]),
                                            .B(encode_v[249])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v250 (
                                            .F(comp_v[250]),
                                            .B(encode_v[250])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v251 (
                                            .F(comp_v[251]),
                                            .B(encode_v[251])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v252 (
                                            .F(comp_v[252]),
                                            .B(encode_v[252])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v253 (
                                            .F(comp_v[253]),
                                            .B(encode_v[253])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v254 (
                                            .F(comp_v[254]),
                                            .B(encode_v[254])
                                        );
                                        
                                        encode #(.D(4),.BYTE_LEN(32))enc_v255 (
                                            .F(comp_v[255]),
                                            .B(encode_v[255])
                                        );
always_ff @(posedge clk or posedge rst) begin
                                     if (rst) begin
                                     ntt_started <=0;
                                         all_shake_done <= 0;
                                         mul <= 0;
                          //                       start_encode <= 0;
                                                 start_parse  <= 0;
                                                 start_cbd    <= 0;
                                                 start_prf    <= 0;
                          //                       start_ntt <= 0;
                                     end else begin
                          //           start_mul <=0;
                          //           start_encode<=0;
                          //ntt_started <=0;
//                          start_ntt <= 0;
                          
//                                     start_mul    <= 0;
                          //                   start_encode <= 0;
                                             start_parse  <= 0;
                                             start_cbd    <= 0;
                                             start_prf    <= 0;
                                      start1 <= 1;
                                     zetas[0] = 17; zetas[1] = 2761; zetas[2] = 583; zetas[3] = 2649; zetas[4] = 1637; zetas[5] = 723; zetas[6] = 2288; zetas[7] = 1100;
                                             zetas[8] = 1409; zetas[9] = 2662; zetas[10] = 3281; zetas[11] = 233; zetas[12] = 756; zetas[13] = 2156; zetas[14] = 3015; zetas[15] = 3050;
                                             zetas[16] = 1703; zetas[17] = 1651; zetas[18] = 2789; zetas[19] = 1789; zetas[20] = 1847; zetas[21] = 952; zetas[22] = 1461; zetas[23] = 2687;
                                             zetas[24] = 939; zetas[25] = 2308; zetas[26] = 2437; zetas[27] = 2388; zetas[28] = 733; zetas[29] = 2337; zetas[30] = 268; zetas[31] = 641;
                                             zetas[32] = 1584; zetas[33] = 2298; zetas[34] = 2037; zetas[35] = 3220; zetas[36] = 375; zetas[37] = 2549; zetas[38] = 2090; zetas[39] = 1645;
                                             zetas[40] = 1063; zetas[41] = 319; zetas[42] = 2773; zetas[43] = 757; zetas[44] = 2099; zetas[45] = 561; zetas[46] = 2466; zetas[47] = 2594;
                                             zetas[48] = 2804; zetas[49] = 1092; zetas[50] = 403; zetas[51] = 1026; zetas[52] = 1143; zetas[53] = 2150; zetas[54] = 2775; zetas[55] = 886;
                                             zetas[56] = 1722; zetas[57] = 1212; zetas[58] = 1874; zetas[59] = 1029; zetas[60] = 2110; zetas[61] = 2935; zetas[62] = 885; zetas[63] = 2154;
                                             zetas[64] = 289; zetas[65] = 331; zetas[66] = 3253; zetas[67] = 1756; zetas[68] = 1197; zetas[69] = 2304; zetas[70] = 2277; zetas[71] = 2055;
                                             zetas[72] = 650; zetas[73] = 1977; zetas[74] = 2513; zetas[75] = 632; zetas[76] = 2865; zetas[77] = 33; zetas[78] = 1320; zetas[79] = 1915;
                                             zetas[80] = 2319; zetas[81] = 1435; zetas[82] = 807; zetas[83] = 452; zetas[84] = 1438; zetas[85] = 2868; zetas[86] = 1534; zetas[87] = 2402;
                                             zetas[88] = 2647; zetas[89] = 2617; zetas[90] = 1481; zetas[91] = 648; zetas[92] = 2474; zetas[93] = 3110; zetas[94] = 1227; zetas[95] = 910;
                                             zetas[96] = 296; zetas[97] = 2447; zetas[98] = 1339; zetas[99] = 1476; zetas[100] = 3046; zetas[101] = 56; zetas[102] = 2240; zetas[103] = 1333;
                                             zetas[104] = 1426; zetas[105] = 2094; zetas[106] = 535; zetas[107] = 2882; zetas[108] = 2393; zetas[109] = 2879; zetas[110] = 1974; zetas[111] = 821;
                                             zetas[112] = 1062; zetas[113] = 1919; zetas[114] = 193; zetas[115] = 797; zetas[116] = 2786; zetas[117] = 3260; zetas[118] = 569; zetas[119] = 1746;
                                             zetas[120] = 2642; zetas[121] = 630; zetas[122] = 1897; zetas[123] = 848; zetas[124] = 2580; zetas[125] = 3289; zetas[126] = 1729; zetas[127] = 3328;
                                      zetas[17] = 2637;
                                   
                                   
                                    for (int i = 0; i < 768; i = i + 1) begin
                                                     
                                                                    parse_array1[i] = xof[(i+1)*8-1 -: 8];
                                                                     parse_array2[i] = xof2[(i+1)*8-1 -: 8];
                                                                      parse_array3[i] = xof3[(i+1)*8-1 -: 8];
                                                                       parse_array4[i] = xof4[(i+1)*8-1 -: 8];
                                                                        parse_array5[i] = xof5[(i+1)*8-1 -: 8];
                                                                         parse_array6[i] = xof6[(i+1)*8-1 -: 8];
                                                                          parse_array7[i] = xof7[(i+1)*8-1 -: 8];
                                                                           parse_array8[i] = xof8[(i+1)*8-1 -: 8];
                                                                            parse_array9[i] = xof9[(i+1)*8-1 -: 8];
                                                                       
                                     end
                                      if (done0_shake && done1_shake && done2_shake && done3_shake
                                                       && done6_shake && done7_shake && done8_shake  ) begin
                                                       start_parse <= 1;
                                                       start1 <= 0; 
                                                   end
                                                   
                                      if (done0 && done1 && done2 && done3 && done4 && done5 && done6 && done7 && done8 && !done9_shake && !done10_shake && !done11_shake && !done12_shake && !done13_shake && !done14_shake) begin
                                                                                start_parse <= 0;
                                                                                start_prf <= 1;
                                                                                 
                                                                            end
                            for (int i = 0; i < 128; i++) begin
                                                       prf_bytes_0[i] = prf_0[8*i +: 8];
                                                       prf_bytes_1[i] = prf_1[8*i +: 8];
                                                       prf_bytes_2[i] = prf_2[8*i +: 8];
                                                       prf_bytes_3[i] = prf_3[8*i +: 8];
                                                       prf_bytes_4[i] = prf_4[8*i +: 8];
                                                       prf_bytes_5[i] = prf_5[8*i +: 8];
                                                       prf_bytes_6[i] = prf_6[8*i +: 8];
                                                   end
                          //            
                                            if (done0_shake && done1_shake && done2_shake && done3_shake &&
                                                done4_shake && done5_shake && done6_shake && done7_shake && done8_shake) begin
                                                all_shake_done <= 1;
                                                start1 <= 0; 
                                            end else begin
                                                all_shake_done <= 0; 
                                            end
                                       
                                             if (done0_mul && done1_mul && done2_mul && done3_mul && done4_mul && done5_mul && done6_mul && done7_mul && done8_mul) begin
                                                                                                                                           mul_add[0][0] <= ((mult_out_00[0] + mult_out_01[0] + mult_out_02[0])%3329);
                                                                                                                                           mul_add[0][1] <= ((mult_out_00[1] + mult_out_01[1] + mult_out_02[1])%3329) ;
                                                                                                                                           mul_add[0][2] <= ((mult_out_00[2] + mult_out_01[2] + mult_out_02[2])%3329) ;
                                                                                                                                           mul_add[0][3] <= ((mult_out_00[3] + mult_out_01[3] + mult_out_02[3])%3329) ;
                                                                                                                                           mul_add[0][4] <= ((mult_out_00[4] + mult_out_01[4] + mult_out_02[4])%3329) ;
                                                                                                                                           mul_add[0][5]<=((mult_out_00[5] + mult_out_01[5] + mult_out_02[5])%3329) ;
                                                                                                                                           mul_add[0][6]<=((mult_out_00[6] + mult_out_01[6] + mult_out_02[6])%3329);
                                                                                                                                           mul_add[0][7]<=((mult_out_00[7] + mult_out_01[7] + mult_out_02[7])%3329) ;
                                                                                                                                           mul_add[0][8]<=((mult_out_00[8] + mult_out_01[8] + mult_out_02[8])%3329);
                                                                                                                                           mul_add[0][9]<=((mult_out_00[9] + mult_out_01[9] + mult_out_02[9])%3329) ;
                                                                                                                                           mul_add[0][10]<=((mult_out_00[10] + mult_out_01[10] + mult_out_02[10])%3329) ;
                                                                                                                                           mul_add[0][11]<=((mult_out_00[11] + mult_out_01[11] + mult_out_02[11])%3329) ;
                                                                                                                                           mul_add[0][12]<=((mult_out_00[12] + mult_out_01[12] + mult_out_02[12])%3329) ;
                                                                                                                                           mul_add[0][13]<=((mult_out_00[13] + mult_out_01[13] + mult_out_02[13])%3329) ;
                                                                                                                                           mul_add[0][14]<=((mult_out_00[14] + mult_out_01[14] + mult_out_02[14])%3329) ;
                                                                                                                                           mul_add[0][15]<=((mult_out_00[15] + mult_out_01[15] + mult_out_02[15])%3329) ;
                                                                                                                                           mul_add[0][16]<=((mult_out_00[16] + mult_out_01[16] + mult_out_02[16])%3329) ;
                                                                                                                                           mul_add[0][17]<=((mult_out_00[17] + mult_out_01[17] + mult_out_02[17])%3329) ;
                                                                                                                                           mul_add[0][18]<=((mult_out_00[18] + mult_out_01[18] + mult_out_02[18])%3329) ;
                                                                                                                                           mul_add[0][19]<=((mult_out_00[19] + mult_out_01[19] + mult_out_02[19])%3329) ;
                                                                                                                                           mul_add[0][20]<=((mult_out_00[20] + mult_out_01[20] + mult_out_02[20])%3329) ;
                                                                                                                                           mul_add[0][21]<=((mult_out_00[21] + mult_out_01[21] + mult_out_02[21])%3329) ;
                                                                                                                                           mul_add[0][22]<=((mult_out_00[22] + mult_out_01[22] + mult_out_02[22])%3329) ;
                                                                                                                                           mul_add[0][23]<=((mult_out_00[23] + mult_out_01[23] + mult_out_02[23])%3329) ;
                                                                                                                                           mul_add[0][24]<=((mult_out_00[24] + mult_out_01[24] + mult_out_02[24])%3329) ;
                                                                                                                                           mul_add[0][25]<=((mult_out_00[25] + mult_out_01[25] + mult_out_02[25])%3329) ;
                                                                                                                                           mul_add[0][26]<=((mult_out_00[26] + mult_out_01[26] + mult_out_02[26])%3329) ;
                                                                                                                                           mul_add[0][27]<=((mult_out_00[27] + mult_out_01[27] + mult_out_02[27])%3329) ;
                                                                                                                                           mul_add[0][28]<=((mult_out_00[28] + mult_out_01[28] + mult_out_02[28])%3329) ;
                                                                                                                                           mul_add[0][29]<=((mult_out_00[29] + mult_out_01[29] + mult_out_02[29])%3329) ;
                                                                                                                                           mul_add[0][30]<=((mult_out_00[30] + mult_out_01[30] + mult_out_02[30])%3329) ;
                                                                                                                                           mul_add[0][31]<=((mult_out_00[31] + mult_out_01[31] + mult_out_02[31])%3329) ;
                                                                                                                                           mul_add[0][32]<=((mult_out_00[32] + mult_out_01[32] + mult_out_02[32])%3329) ;
                                                                                                                                           mul_add[0][33]<=((mult_out_00[33] + mult_out_01[33] + mult_out_02[33])%3329) ;
                                                                                                                                           mul_add[0][34]<=((mult_out_00[34] + mult_out_01[34] + mult_out_02[34])%3329) ;
                                                                                                                                           mul_add[0][35]<=((mult_out_00[35] + mult_out_01[35] + mult_out_02[35])%3329) ;
                                                                                                                                           mul_add[0][36]<=((mult_out_00[36] + mult_out_01[36] + mult_out_02[36])%3329) ;
                                                                                                                                           mul_add[0][37]<=((mult_out_00[37] + mult_out_01[37] + mult_out_02[37])%3329) ;
                                                                                                                                           mul_add[0][38]<=((mult_out_00[38] + mult_out_01[38] + mult_out_02[38])%3329) ;
                                                                                                                                           mul_add[0][39]<=((mult_out_00[39] + mult_out_01[39] + mult_out_02[39])%3329) ;
                                                                                                                                           mul_add[0][40]<=((mult_out_00[40] + mult_out_01[40] + mult_out_02[40])%3329) ;
                                                                                                                                           mul_add[0][41]<=((mult_out_00[41] + mult_out_01[41] + mult_out_02[41])%3329) ;
                                                                                                                                           mul_add[0][42]<=((mult_out_00[42] + mult_out_01[42] + mult_out_02[42])%3329) ;
                                                                                                                                           mul_add[0][43]<=((mult_out_00[43] + mult_out_01[43] + mult_out_02[43])%3329) ;
                                                                                                                                           mul_add[0][44]<=((mult_out_00[44] + mult_out_01[44] + mult_out_02[44])%3329) ;
                                                                                                                                           mul_add[0][45]<=((mult_out_00[45] + mult_out_01[45] + mult_out_02[45])%3329) ;
                                                                                                                                           mul_add[0][46]<=((mult_out_00[46] + mult_out_01[46] + mult_out_02[46])%3329) ;
                                                                                                                                           mul_add[0][47]<=((mult_out_00[47] + mult_out_01[47] + mult_out_02[47])%3329) ;
                                                                                                                                           mul_add[0][48]<=((mult_out_00[48] + mult_out_01[48] + mult_out_02[48])%3329) ;
                                                                                                                                           mul_add[0][49]<=((mult_out_00[49] + mult_out_01[49] + mult_out_02[49])%3329) ;
                                                                                                                                           mul_add[0][50]<=((mult_out_00[50] + mult_out_01[50] + mult_out_02[50])%3329) ;
                                                                                                                                           mul_add[0][51]<=((mult_out_00[51] + mult_out_01[51] + mult_out_02[51])%3329) ;
                                                                                                                                           mul_add[0][52]<=((mult_out_00[52] + mult_out_01[52] + mult_out_02[52])%3329) ;
                                                                                                                                           mul_add[0][53]<=((mult_out_00[53] + mult_out_01[53] + mult_out_02[53])%3329) ;
                                                                                                                                           mul_add[0][54]<=((mult_out_00[54] + mult_out_01[54] + mult_out_02[54])%3329) ;
                                                                                                                                           mul_add[0][55]<=((mult_out_00[55] + mult_out_01[55] + mult_out_02[55])%3329) ;
                                                                                                                                           mul_add[0][56]<=((mult_out_00[56] + mult_out_01[56] + mult_out_02[56])%3329) ;
                                                                                                                                           mul_add[0][57]<=((mult_out_00[57] + mult_out_01[57] + mult_out_02[57])%3329) ;
                                                                                                                                           mul_add[0][58]<=((mult_out_00[58] + mult_out_01[58] + mult_out_02[58])%3329) ;
                                                                                                                                           mul_add[0][59]<=((mult_out_00[59] + mult_out_01[59] + mult_out_02[59])%3329) ;
                                                                                                                                           mul_add[0][60]<=((mult_out_00[60] + mult_out_01[60] + mult_out_02[60])%3329) ;
                                                                                                                                           mul_add[0][61]<=((mult_out_00[61] + mult_out_01[61] + mult_out_02[61])%3329) ;
                                                                                                                                           mul_add[0][62]<=((mult_out_00[62] + mult_out_01[62] + mult_out_02[62])%3329) ;
                                                                                                                                           mul_add[0][63]<=((mult_out_00[63] + mult_out_01[63] + mult_out_02[63])%3329) ;
                                                                                                                                           mul_add[0][64]<=((mult_out_00[64] + mult_out_01[64] + mult_out_02[64])%3329) ;
                                                                                                                                           mul_add[0][65]<=((mult_out_00[65] + mult_out_01[65] + mult_out_02[65])%3329) ;
                                                                                                                                           mul_add[0][66]<=((mult_out_00[66] + mult_out_01[66] + mult_out_02[66])%3329) ;
                                                                                                                                           mul_add[0][67]<=((mult_out_00[67] + mult_out_01[67] + mult_out_02[67])%3329) ;
                                                                                                                                           mul_add[0][68]<=((mult_out_00[68] + mult_out_01[68] + mult_out_02[68])%3329) ;
                                                                                                                                           mul_add[0][69]<=((mult_out_00[69] + mult_out_01[69] + mult_out_02[69])%3329) ;
                                                                                                                                           mul_add[0][70]<=((mult_out_00[70] + mult_out_01[70] + mult_out_02[70])%3329) ;
                                                                                                                                           mul_add[0][71]<=((mult_out_00[71] + mult_out_01[71] + mult_out_02[71])%3329) ;
                                                                                                                                           mul_add[0][72]<=((mult_out_00[72] + mult_out_01[72] + mult_out_02[72])%3329) ;
                                                                                                                                           mul_add[0][73]<=((mult_out_00[73] + mult_out_01[73] + mult_out_02[73])%3329) ;
                                                                                                                                           mul_add[0][74]<=((mult_out_00[74] + mult_out_01[74] + mult_out_02[74])%3329) ;
                                                                                                                                           mul_add[0][75]<=((mult_out_00[75] + mult_out_01[75] + mult_out_02[75])%3329) ;
                                                                                                                                           mul_add[0][76]<=((mult_out_00[76] + mult_out_01[76] + mult_out_02[76])%3329) ;
                                                                                                                                           mul_add[0][77]<=((mult_out_00[77] + mult_out_01[77] + mult_out_02[77])%3329) ;
                                                                                                                                           mul_add[0][78]<=((mult_out_00[78] + mult_out_01[78] + mult_out_02[78])%3329) ;
                                                                                                                                           mul_add[0][79]<=((mult_out_00[79] + mult_out_01[79] + mult_out_02[79])%3329) ;
                                                                                                                                           mul_add[0][80]<=((mult_out_00[80] + mult_out_01[80] + mult_out_02[80])%3329) ;
                                                                                                                                           mul_add[0][81]<=((mult_out_00[81] + mult_out_01[81] + mult_out_02[81])%3329) ;
                                                                                                                                           mul_add[0][82]<=((mult_out_00[82] + mult_out_01[82] + mult_out_02[82])%3329) ;
                                                                                                                                           mul_add[0][83]<=((mult_out_00[83] + mult_out_01[83] + mult_out_02[83])%3329) ;
                                                                                                                                           mul_add[0][84]<=((mult_out_00[84] + mult_out_01[84] + mult_out_02[84])%3329) ;
                                                                                                                                           mul_add[0][85]<=((mult_out_00[85] + mult_out_01[85] + mult_out_02[85])%3329) ;
                                                                                                                                           mul_add[0][86]<=((mult_out_00[86] + mult_out_01[86] + mult_out_02[86])%3329) ;
                                                                                                                                           mul_add[0][87]<=((mult_out_00[87] + mult_out_01[87] + mult_out_02[87])%3329) ;
                                                                                                                                           mul_add[0][88]<=((mult_out_00[88] + mult_out_01[88] + mult_out_02[88])%3329) ;
                                                                                                                                           mul_add[0][89]<=((mult_out_00[89] + mult_out_01[89] + mult_out_02[89])%3329) ;
                                                                                                                                           mul_add[0][90]<=((mult_out_00[90] + mult_out_01[90] + mult_out_02[90])%3329) ;
                                                                                                                                           mul_add[0][91]<=((mult_out_00[91] + mult_out_01[91] + mult_out_02[91])%3329) ;
                                                                                                                                           mul_add[0][92]<=((mult_out_00[92] + mult_out_01[92] + mult_out_02[92])%3329) ;
                                                                                                                                           mul_add[0][93]<=((mult_out_00[93] + mult_out_01[93] + mult_out_02[93])%3329) ;
                                                                                                                                           mul_add[0][94]<=((mult_out_00[94] + mult_out_01[94] + mult_out_02[94])%3329) ;
                                                                                                                                           mul_add[0][95]<=((mult_out_00[95] + mult_out_01[95] + mult_out_02[95])%3329) ;
                                                                                                                                           mul_add[0][96]<=((mult_out_00[96] + mult_out_01[96] + mult_out_02[96])%3329) ;
                                                                                                                                           mul_add[0][97]<=((mult_out_00[97] + mult_out_01[97] + mult_out_02[97])%3329) ;
                                                                                                                                           mul_add[0][98]<=((mult_out_00[98] + mult_out_01[98] + mult_out_02[98])%3329) ;
                                                                                                                                           mul_add[0][99]<=((mult_out_00[99] + mult_out_01[99] + mult_out_02[99])%3329) ;
                                                                                                                                           mul_add[0][100]<=((mult_out_00[100] + mult_out_01[100] + mult_out_02[100])%3329) ;
                                                                                                                                           mul_add[0][101]<=((mult_out_00[101] + mult_out_01[101] + mult_out_02[101])%3329) ;
                                                                                                                                           mul_add[0][102]<=((mult_out_00[102] + mult_out_01[102] + mult_out_02[102])%3329) ;
                                                                                                                                           mul_add[0][103]<=((mult_out_00[103] + mult_out_01[103] + mult_out_02[103])%3329) ;
                                                                                                                                           mul_add[0][104]<=((mult_out_00[104] + mult_out_01[104] + mult_out_02[104])%3329) ;
                                                                                                                                           mul_add[0][105]<=((mult_out_00[105] + mult_out_01[105] + mult_out_02[105])%3329) ;
                                                                                                                                           mul_add[0][106]<=((mult_out_00[106] + mult_out_01[106] + mult_out_02[106])%3329) ;
                                                                                                                                           mul_add[0][107]<=((mult_out_00[107] + mult_out_01[107] + mult_out_02[107])%3329) ;
                                                                                                                                           mul_add[0][108]<=((mult_out_00[108] + mult_out_01[108] + mult_out_02[108])%3329) ;
                                                                                                                                           mul_add[0][109]<=((mult_out_00[109] + mult_out_01[109] + mult_out_02[109])%3329) ;
                                                                                                                                           mul_add[0][110]<=((mult_out_00[110] + mult_out_01[110] + mult_out_02[110])%3329) ;
                                                                                                                                           mul_add[0][111]<=((mult_out_00[111] + mult_out_01[111] + mult_out_02[111])%3329) ;
                                                                                                                                           mul_add[0][112]<=((mult_out_00[112] + mult_out_01[112] + mult_out_02[112])%3329) ;
                                                                                                                                           mul_add[0][113]<=((mult_out_00[113] + mult_out_01[113] + mult_out_02[113])%3329) ;
                                                                                                                                           mul_add[0][114]<=((mult_out_00[114] + mult_out_01[114] + mult_out_02[114])%3329) ;
                                                                                                                                           mul_add[0][115]<=((mult_out_00[115] + mult_out_01[115] + mult_out_02[115])%3329) ;
                                                                                                                                           mul_add[0][116]<=((mult_out_00[116] + mult_out_01[116] + mult_out_02[116])%3329) ;
                                                                                                                                           mul_add[0][117]<=((mult_out_00[117] + mult_out_01[117] + mult_out_02[117])%3329) ;
                                                                                                                                           mul_add[0][118]<=((mult_out_00[118] + mult_out_01[118] + mult_out_02[118])%3329) ;
                                                                                                                                           mul_add[0][119]<=((mult_out_00[119] + mult_out_01[119] + mult_out_02[119])%3329) ;
                                                                                                                                           mul_add[0][120]<=((mult_out_00[120] + mult_out_01[120] + mult_out_02[120])%3329) ;
                                                                                                                                           mul_add[0][121]<=((mult_out_00[121] + mult_out_01[121] + mult_out_02[121])%3329) ;
                                                                                                                                           mul_add[0][122]<=((mult_out_00[122] + mult_out_01[122] + mult_out_02[122])%3329) ;
                                                                                                                                           mul_add[0][123]<=((mult_out_00[123] + mult_out_01[123] + mult_out_02[123])%3329) ;
                                                                                                                                           mul_add[0][124]<=((mult_out_00[124] + mult_out_01[124] + mult_out_02[124])%3329) ;
                                                                                                                                           mul_add[0][125]<=((mult_out_00[125] + mult_out_01[125] + mult_out_02[125])%3329) ;
                                                                                                                                           mul_add[0][126]<=((mult_out_00[126] + mult_out_01[126] + mult_out_02[126])%3329) ;
                                                                                                                                           mul_add[0][127]<=((mult_out_00[127] + mult_out_01[127] + mult_out_02[127])%3329) ;
                                                                                                                                           mul_add[0][128]<=((mult_out_00[128] + mult_out_01[128] + mult_out_02[128])%3329) ;
                                                                                                                                           mul_add[0][129]<=((mult_out_00[129] + mult_out_01[129] + mult_out_02[129])%3329) ;
                                                                                                                                           mul_add[0][130]<=((mult_out_00[130] + mult_out_01[130] + mult_out_02[130])%3329) ;
                                                                                                                                           mul_add[0][131]<=((mult_out_00[131] + mult_out_01[131] + mult_out_02[131])%3329) ;
                                                                                                                                           mul_add[0][132]<=((mult_out_00[132] + mult_out_01[132] + mult_out_02[132])%3329) ;
                                                                                                                                           mul_add[0][133]<=((mult_out_00[133] + mult_out_01[133] + mult_out_02[133])%3329) ;
                                                                                                                                           mul_add[0][134]<=((mult_out_00[134] + mult_out_01[134] + mult_out_02[134])%3329) ;
                                                                                                                                           mul_add[0][135]<=((mult_out_00[135] + mult_out_01[135] + mult_out_02[135])%3329) ;
                                                                                                                                           mul_add[0][136]<=((mult_out_00[136] + mult_out_01[136] + mult_out_02[136])%3329) ;
                                                                                                                                           mul_add[0][137]<=((mult_out_00[137] + mult_out_01[137] + mult_out_02[137])%3329) ;
                                                                                                                                           mul_add[0][138]<=((mult_out_00[138] + mult_out_01[138] + mult_out_02[138])%3329) ;
                                                                                                                                           mul_add[0][139]<=((mult_out_00[139] + mult_out_01[139] + mult_out_02[139])%3329) ;
                                                                                                                                           mul_add[0][140]<=((mult_out_00[140] + mult_out_01[140] + mult_out_02[140])%3329) ;
                                                                                                                                           mul_add[0][141]<=((mult_out_00[141] + mult_out_01[141] + mult_out_02[141])%3329) ;
                                                                                                                                           mul_add[0][142]<=((mult_out_00[142] + mult_out_01[142] + mult_out_02[142])%3329) ;
                                                                                                                                           mul_add[0][143]<=((mult_out_00[143] + mult_out_01[143] + mult_out_02[143])%3329) ;
                                                                                                                                           mul_add[0][144]<=((mult_out_00[144] + mult_out_01[144] + mult_out_02[144])%3329) ;
                                                                                                                                           mul_add[0][145]<=((mult_out_00[145] + mult_out_01[145] + mult_out_02[145])%3329) ;
                                                                                                                                           mul_add[0][146]<=((mult_out_00[146] + mult_out_01[146] + mult_out_02[146])%3329) ;
                                                                                                                                           mul_add[0][147]<=((mult_out_00[147] + mult_out_01[147] + mult_out_02[147])%3329) ;
                                                                                                                                           mul_add[0][148]<=((mult_out_00[148] + mult_out_01[148] + mult_out_02[148])%3329) ;
                                                                                                                                           mul_add[0][149]<=((mult_out_00[149] + mult_out_01[149] + mult_out_02[149])%3329) ;
                                                                                                                                           mul_add[0][150]<=((mult_out_00[150] + mult_out_01[150] + mult_out_02[150])%3329) ;
                                                                                                                                           mul_add[0][151]<=((mult_out_00[151] + mult_out_01[151] + mult_out_02[151])%3329) ;
                                                                                                                                           mul_add[0][152]<=((mult_out_00[152] + mult_out_01[152] + mult_out_02[152])%3329) ;
                                                                                                                                           mul_add[0][153]<=((mult_out_00[153] + mult_out_01[153] + mult_out_02[153])%3329) ;
                                                                                                                                           mul_add[0][154]<=((mult_out_00[154] + mult_out_01[154] + mult_out_02[154])%3329) ;
                                                                                                                                           mul_add[0][155]<=((mult_out_00[155] + mult_out_01[155] + mult_out_02[155])%3329) ;
                                                                                                                                           mul_add[0][156]<=((mult_out_00[156] + mult_out_01[156] + mult_out_02[156])%3329) ;
                                                                                                                                           mul_add[0][157]<=((mult_out_00[157] + mult_out_01[157] + mult_out_02[157])%3329) ;
                                                                                                                                           mul_add[0][158]<=((mult_out_00[158] + mult_out_01[158] + mult_out_02[158])%3329) ;
                                                                                                                                           mul_add[0][159]<=((mult_out_00[159] + mult_out_01[159] + mult_out_02[159])%3329) ;
                                                                                                                                           mul_add[0][160]<=((mult_out_00[160] + mult_out_01[160] + mult_out_02[160])%3329) ;
                                                                                                                                           mul_add[0][161]<=((mult_out_00[161] + mult_out_01[161] + mult_out_02[161])%3329) ;
                                                                                                                                           mul_add[0][162]<=((mult_out_00[162] + mult_out_01[162] + mult_out_02[162])%3329) ;
                                                                                                                                           mul_add[0][163]<=((mult_out_00[163] + mult_out_01[163] + mult_out_02[163])%3329) ;
                                                                                                                                           mul_add[0][164]<=((mult_out_00[164] + mult_out_01[164] + mult_out_02[164])%3329) ;
                                                                                                                                           mul_add[0][165]<=((mult_out_00[165] + mult_out_01[165] + mult_out_02[165])%3329) ;
                                                                                                                                           mul_add[0][166]<=((mult_out_00[166] + mult_out_01[166] + mult_out_02[166])%3329) ;
                                                                                                                                           mul_add[0][167]<=((mult_out_00[167] + mult_out_01[167] + mult_out_02[167])%3329) ;
                                                                                                                                           mul_add[0][168]<=((mult_out_00[168] + mult_out_01[168] + mult_out_02[168])%3329) ;
                                                                                                                                           mul_add[0][169]<=((mult_out_00[169] + mult_out_01[169] + mult_out_02[169])%3329) ;
                                                                                                                                           mul_add[0][170]<=((mult_out_00[170] + mult_out_01[170] + mult_out_02[170])%3329) ;
                                                                                                                                           mul_add[0][171]<=((mult_out_00[171] + mult_out_01[171] + mult_out_02[171])%3329) ;
                                                                                                                                           mul_add[0][172]<=((mult_out_00[172] + mult_out_01[172] + mult_out_02[172])%3329) ;
                                                                                                                                           mul_add[0][173]<=((mult_out_00[173] + mult_out_01[173] + mult_out_02[173])%3329) ;
                                                                                                                                           mul_add[0][174]<=((mult_out_00[174] + mult_out_01[174] + mult_out_02[174])%3329) ;
                                                                                                                                           mul_add[0][175]<=((mult_out_00[175] + mult_out_01[175] + mult_out_02[175])%3329) ;
                                                                                                                                           mul_add[0][176]<=((mult_out_00[176] + mult_out_01[176] + mult_out_02[176])%3329) ;
                                                                                                                                           mul_add[0][177]<=((mult_out_00[177] + mult_out_01[177] + mult_out_02[177])%3329) ;
                                                                                                                                           mul_add[0][178]<=((mult_out_00[178] + mult_out_01[178] + mult_out_02[178])%3329) ;
                                                                                                                                           mul_add[0][179]<=((mult_out_00[179] + mult_out_01[179] + mult_out_02[179])%3329) ;
                                                                                                                                           mul_add[0][180]<=((mult_out_00[180] + mult_out_01[180] + mult_out_02[180])%3329) ;
                                                                                                                                           mul_add[0][181]<=((mult_out_00[181] + mult_out_01[181] + mult_out_02[181])%3329) ;
                                                                                                                                           mul_add[0][182]<=((mult_out_00[182] + mult_out_01[182] + mult_out_02[182])%3329) ;
                                                                                                                                           mul_add[0][183]<=((mult_out_00[183] + mult_out_01[183] + mult_out_02[183])%3329) ;
                                                                                                                                           mul_add[0][184]<=((mult_out_00[184] + mult_out_01[184] + mult_out_02[184])%3329) ;
                                                                                                                                           mul_add[0][185]<=((mult_out_00[185] + mult_out_01[185] + mult_out_02[185])%3329) ;
                                                                                                                                           mul_add[0][186]<=((mult_out_00[186] + mult_out_01[186] + mult_out_02[186])%3329) ;
                                                                                                                                           mul_add[0][187]<=((mult_out_00[187] + mult_out_01[187] + mult_out_02[187])%3329) ;
                                                                                                                                           mul_add[0][188]<=((mult_out_00[188] + mult_out_01[188] + mult_out_02[188])%3329) ;
                                                                                                                                           mul_add[0][189]<=((mult_out_00[189] + mult_out_01[189] + mult_out_02[189])%3329) ;
                                                                                                                                           mul_add[0][190]<=((mult_out_00[190] + mult_out_01[190] + mult_out_02[190])%3329) ;
                                                                                                                                           mul_add[0][191]<=((mult_out_00[191] + mult_out_01[191] + mult_out_02[191])%3329) ;
                                                                                                                                           mul_add[0][192]<=((mult_out_00[192] + mult_out_01[192] + mult_out_02[192])%3329) ;
                                                                                                                                           mul_add[0][193]<=((mult_out_00[193] + mult_out_01[193] + mult_out_02[193])%3329) ;
                                                                                                                                           mul_add[0][194]<=((mult_out_00[194] + mult_out_01[194] + mult_out_02[194])%3329) ;
                                                                                                                                           mul_add[0][195]<=((mult_out_00[195] + mult_out_01[195] + mult_out_02[195])%3329) ;
                                                                                                                                           mul_add[0][196]<=((mult_out_00[196] + mult_out_01[196] + mult_out_02[196])%3329) ;
                                                                                                                                           mul_add[0][197]<=((mult_out_00[197] + mult_out_01[197] + mult_out_02[197])%3329) ;
                                                                                                                                           mul_add[0][198]<=((mult_out_00[198] + mult_out_01[198] + mult_out_02[198])%3329) ;
                                                                                                                                           mul_add[0][199]<=((mult_out_00[199] + mult_out_01[199] + mult_out_02[199])%3329) ;
                                                                                                                                           mul_add[0][200]<=((mult_out_00[200] + mult_out_01[200] + mult_out_02[200])%3329) ;
                                                                                                                                           mul_add[0][201]<=((mult_out_00[201] + mult_out_01[201] + mult_out_02[201])%3329) ;
                                                                                                                                           mul_add[0][202]<=((mult_out_00[202] + mult_out_01[202] + mult_out_02[202])%3329) ;
                                                                                                                                           mul_add[0][203]<=((mult_out_00[203] + mult_out_01[203] + mult_out_02[203])%3329) ;
                                                                                                                                           mul_add[0][204]<=((mult_out_00[204] + mult_out_01[204] + mult_out_02[204])%3329) ;
                                                                                                                                           mul_add[0][205]<=((mult_out_00[205] + mult_out_01[205] + mult_out_02[205])%3329) ;
                                                                                                                                           mul_add[0][206]<=((mult_out_00[206] + mult_out_01[206] + mult_out_02[206])%3329) ;
                                                                                                                                           mul_add[0][207]<=((mult_out_00[207] + mult_out_01[207] + mult_out_02[207])%3329) ;
                                                                                                                                           mul_add[0][208]<=((mult_out_00[208] + mult_out_01[208] + mult_out_02[208])%3329) ;
                                                                                                                                           mul_add[0][209]<=((mult_out_00[209] + mult_out_01[209] + mult_out_02[209])%3329) ;
                                                                                                                                           mul_add[0][210]<=((mult_out_00[210] + mult_out_01[210] + mult_out_02[210])%3329) ;
                                                                                                                                           mul_add[0][211]<=((mult_out_00[211] + mult_out_01[211] + mult_out_02[211])%3329) ;
                                                                                                                                           mul_add[0][212]<=((mult_out_00[212] + mult_out_01[212] + mult_out_02[212])%3329) ;
                                                                                                                                           mul_add[0][213]<=((mult_out_00[213] + mult_out_01[213] + mult_out_02[213])%3329) ;
                                                                                                                                           mul_add[0][214]<=((mult_out_00[214] + mult_out_01[214] + mult_out_02[214])%3329) ;
                                                                                                                                           mul_add[0][215]<=((mult_out_00[215] + mult_out_01[215] + mult_out_02[215])%3329) ;
                                                                                                                                           mul_add[0][216]<=((mult_out_00[216] + mult_out_01[216] + mult_out_02[216])%3329) ;
                                                                                                                                           mul_add[0][217]<=((mult_out_00[217] + mult_out_01[217] + mult_out_02[217])%3329) ;
                                                                                                                                           mul_add[0][218]<=((mult_out_00[218] + mult_out_01[218] + mult_out_02[218])%3329) ;
                                                                                                                                           mul_add[0][219]<=((mult_out_00[219] + mult_out_01[219] + mult_out_02[219])%3329) ;
                                                                                                                                           mul_add[0][220]<=((mult_out_00[220] + mult_out_01[220] + mult_out_02[220])%3329) ;
                                                                                                                                           mul_add[0][221]<=((mult_out_00[221] + mult_out_01[221] + mult_out_02[221])%3329) ;
                                                                                                                                           mul_add[0][222]<=((mult_out_00[222] + mult_out_01[222] + mult_out_02[222])%3329) ;
                                                                                                                                           mul_add[0][223]<=((mult_out_00[223] + mult_out_01[223] + mult_out_02[223])%3329) ;
                                                                                                                                           mul_add[0][224]<=((mult_out_00[224] + mult_out_01[224] + mult_out_02[224])%3329) ;
                                                                                                                                           mul_add[0][225]<=((mult_out_00[225] + mult_out_01[225] + mult_out_02[225])%3329) ;
                                                                                                                                           mul_add[0][226]<=((mult_out_00[226] + mult_out_01[226] + mult_out_02[226])%3329) ;
                                                                                                                                           mul_add[0][227]<=((mult_out_00[227] + mult_out_01[227] + mult_out_02[227])%3329) ;
                                                                                                                                           mul_add[0][228]<=((mult_out_00[228] + mult_out_01[228] + mult_out_02[228])%3329) ;
                                                                                                                                           mul_add[0][229]<=((mult_out_00[229] + mult_out_01[229] + mult_out_02[229])%3329) ;
                                                                                                                                           mul_add[0][230]<=((mult_out_00[230] + mult_out_01[230] + mult_out_02[230])%3329) ;
                                                                                                                                           mul_add[0][231]<=((mult_out_00[231] + mult_out_01[231] + mult_out_02[231])%3329) ;
                                                                                                                                           mul_add[0][232]<=((mult_out_00[232] + mult_out_01[232] + mult_out_02[232])%3329) ;
                                                                                                                                           mul_add[0][233]<=((mult_out_00[233] + mult_out_01[233] + mult_out_02[233])%3329) ;
                                                                                                                                           mul_add[0][234]<=((mult_out_00[234] + mult_out_01[234] + mult_out_02[234])%3329) ;
                                                                                                                                           mul_add[0][235]<=((mult_out_00[235] + mult_out_01[235] + mult_out_02[235])%3329) ;
                                                                                                                                           mul_add[0][236]<=((mult_out_00[236] + mult_out_01[236] + mult_out_02[236])%3329) ;
                                                                                                                                           mul_add[0][237]<=((mult_out_00[237] + mult_out_01[237] + mult_out_02[237])%3329) ;
                                                                                                                                           mul_add[0][238]<=((mult_out_00[238] + mult_out_01[238] + mult_out_02[238])%3329) ;
                                                                                                                                           mul_add[0][239]<=((mult_out_00[239] + mult_out_01[239] + mult_out_02[239])%3329) ;
                                                                                                                                           mul_add[0][240]<=((mult_out_00[240] + mult_out_01[240] + mult_out_02[240])%3329) ;
                                                                                                                                           mul_add[0][241]<=((mult_out_00[241] + mult_out_01[241] + mult_out_02[241])%3329) ;
                                                                                                                                           mul_add[0][242]<=((mult_out_00[242] + mult_out_01[242] + mult_out_02[242])%3329) ;
                                                                                                                                           mul_add[0][243]<=((mult_out_00[243] + mult_out_01[243] + mult_out_02[243])%3329) ;
                                                                                                                                           mul_add[0][244]<=((mult_out_00[244] + mult_out_01[244] + mult_out_02[244])%3329) ;
                                                                                                                                           mul_add[0][245]<=((mult_out_00[245] + mult_out_01[245] + mult_out_02[245])%3329) ;
                                                                                                                                           mul_add[0][246]<=((mult_out_00[246] + mult_out_01[246] + mult_out_02[246])%3329) ;
                                                                                                                                           mul_add[0][247]<=((mult_out_00[247] + mult_out_01[247] + mult_out_02[247])%3329) ;
                                                                                                                                           mul_add[0][248]<=((mult_out_00[248] + mult_out_01[248] + mult_out_02[248])%3329) ;
                                                                                                                                           mul_add[0][249]<=((mult_out_00[249] + mult_out_01[249] + mult_out_02[249])%3329) ;
                                                                                                                                           mul_add[0][250]<=((mult_out_00[250] + mult_out_01[250] + mult_out_02[250])%3329) ;
                                                                                                                                           mul_add[0][251]<=((mult_out_00[251] + mult_out_01[251] + mult_out_02[251])%3329) ;
                                                                                                                                           mul_add[0][252]<=((mult_out_00[252] + mult_out_01[252] + mult_out_02[252])%3329) ;
                                                                                                                                           mul_add[0][253]<=((mult_out_00[253] + mult_out_01[253] + mult_out_02[253])%3329) ;
                                                                                                                                           mul_add[0][254]<=((mult_out_00[254] + mult_out_01[254] + mult_out_02[254])%3329) ;
                                                                                                                                           mul_add[0][255]<=((mult_out_00[255] + mult_out_01[255] + mult_out_02[255])%3329) ;
                                                                                                                                          
                                                                                                                                           mul_add[1][0]<=((mult_out_10[0] + mult_out_11[0] + mult_out_12[0])%3329) ;
                                                                                                                                           mul_add[1][1]<=((mult_out_10[1] + mult_out_11[1] + mult_out_12[1])%3329) ;
                                                                                                                                           mul_add[1][2]<=((mult_out_10[2] + mult_out_11[2] + mult_out_12[2])%3329) ;
                                                                                                                                           mul_add[1][3]<=((mult_out_10[3] + mult_out_11[3] + mult_out_12[3])%3329) ;
                                                                                                                                           mul_add[1][4]<=((mult_out_10[4] + mult_out_11[4] + mult_out_12[4])%3329) ;
                                                                                                                                           mul_add[1][5]<=((mult_out_10[5] + mult_out_11[5] + mult_out_12[5])%3329) ;
                                                                                                                                           mul_add[1][6]<=((mult_out_10[6] + mult_out_11[6] + mult_out_12[6])%3329) ;
                                                                                                                                           mul_add[1][7]<=((mult_out_10[7] + mult_out_11[7] + mult_out_12[7])%3329) ;
                                                                                                                                           mul_add[1][8]<=((mult_out_10[8] + mult_out_11[8] + mult_out_12[8])%3329) ;
                                                                                                                                           mul_add[1][9]<=((mult_out_10[9] + mult_out_11[9] + mult_out_12[9])%3329) ;
                                                                                                                                           mul_add[1][10]<=((mult_out_10[10] + mult_out_11[10] + mult_out_12[10])%3329) ;
                                                                                                                                           mul_add[1][11]<=((mult_out_10[11] + mult_out_11[11] + mult_out_12[11])%3329) ;
                                                                                                                                           mul_add[1][12]<=((mult_out_10[12] + mult_out_11[12] + mult_out_12[12])%3329) ;
                                                                                                                                           mul_add[1][13]<=((mult_out_10[13] + mult_out_11[13] + mult_out_12[13])%3329) ;
                                                                                                                                           mul_add[1][14]<=((mult_out_10[14] + mult_out_11[14] + mult_out_12[14])%3329) ;
                                                                                                                                           mul_add[1][15]<=((mult_out_10[15] + mult_out_11[15] + mult_out_12[15])%3329) ;
                                                                                                                                           mul_add[1][16]<=((mult_out_10[16] + mult_out_11[16] + mult_out_12[16])%3329) ;
                                                                                                                                           mul_add[1][17]<=((mult_out_10[17] + mult_out_11[17] + mult_out_12[17])%3329) ;
                                                                                                                                           mul_add[1][18]<=((mult_out_10[18] + mult_out_11[18] + mult_out_12[18])%3329) ;
                                                                                                                                           mul_add[1][19]<=((mult_out_10[19] + mult_out_11[19] + mult_out_12[19])%3329) ;
                                                                                                                                           mul_add[1][20]<=((mult_out_10[20] + mult_out_11[20] + mult_out_12[20])%3329) ;
                                                                                                                                           mul_add[1][21]<=((mult_out_10[21] + mult_out_11[21] + mult_out_12[21])%3329) ;
                                                                                                                                           mul_add[1][22]<=((mult_out_10[22] + mult_out_11[22] + mult_out_12[22])%3329) ;
                                                                                                                                           mul_add[1][23]<=((mult_out_10[23] + mult_out_11[23] + mult_out_12[23])%3329) ;
                                                                                                                                           mul_add[1][24]<=((mult_out_10[24] + mult_out_11[24] + mult_out_12[24])%3329) ;
                                                                                                                                           mul_add[1][25]<=((mult_out_10[25] + mult_out_11[25] + mult_out_12[25])%3329) ;
                                                                                                                                           mul_add[1][26]<=((mult_out_10[26] + mult_out_11[26] + mult_out_12[26])%3329) ;
                                                                                                                                           mul_add[1][27]<=((mult_out_10[27] + mult_out_11[27] + mult_out_12[27])%3329) ;
                                                                                                                                           mul_add[1][28]<=((mult_out_10[28] + mult_out_11[28] + mult_out_12[28])%3329) ;
                                                                                                                                           mul_add[1][29]<=((mult_out_10[29] + mult_out_11[29] + mult_out_12[29])%3329) ;
                                                                                                                                           mul_add[1][30]<=((mult_out_10[30] + mult_out_11[30] + mult_out_12[30])%3329) ;
                                                                                                                                           mul_add[1][31]<=((mult_out_10[31] + mult_out_11[31] + mult_out_12[31])%3329) ;
                                                                                                                                           mul_add[1][32]<=((mult_out_10[32] + mult_out_11[32] + mult_out_12[32])%3329) ;
                                                                                                                                           mul_add[1][33]<=((mult_out_10[33] + mult_out_11[33] + mult_out_12[33])%3329) ;
                                                                                                                                           mul_add[1][34]<=((mult_out_10[34] + mult_out_11[34] + mult_out_12[34])%3329) ;
                                                                                                                                           mul_add[1][35]<=((mult_out_10[35] + mult_out_11[35] + mult_out_12[35])%3329) ;
                                                                                                                                           mul_add[1][36]<=((mult_out_10[36] + mult_out_11[36] + mult_out_12[36])%3329) ;
                                                                                                                                           mul_add[1][37]<=((mult_out_10[37] + mult_out_11[37] + mult_out_12[37])%3329) ;
                                                                                                                                           mul_add[1][38]<=((mult_out_10[38] + mult_out_11[38] + mult_out_12[38])%3329) ;
                                                                                                                                           mul_add[1][39]<=((mult_out_10[39] + mult_out_11[39] + mult_out_12[39])%3329) ;
                                                                                                                                           mul_add[1][40]<=((mult_out_10[40] + mult_out_11[40] + mult_out_12[40])%3329) ;
                                                                                                                                           mul_add[1][41]<=((mult_out_10[41] + mult_out_11[41] + mult_out_12[41])%3329) ;
                                                                                                                                           mul_add[1][42]<=((mult_out_10[42] + mult_out_11[42] + mult_out_12[42])%3329) ;
                                                                                                                                           mul_add[1][43]<=((mult_out_10[43] + mult_out_11[43] + mult_out_12[43])%3329) ;
                                                                                                                                           mul_add[1][44]<=((mult_out_10[44] + mult_out_11[44] + mult_out_12[44])%3329) ;
                                                                                                                                           mul_add[1][45]<=((mult_out_10[45] + mult_out_11[45] + mult_out_12[45])%3329) ;
                                                                                                                                           mul_add[1][46]<=((mult_out_10[46] + mult_out_11[46] + mult_out_12[46])%3329) ;
                                                                                                                                           mul_add[1][47]<=((mult_out_10[47] + mult_out_11[47] + mult_out_12[47])%3329) ;
                                                                                                                                           mul_add[1][48]<=((mult_out_10[48] + mult_out_11[48] + mult_out_12[48])%3329) ;
                                                                                                                                           mul_add[1][49]<=((mult_out_10[49] + mult_out_11[49] + mult_out_12[49])%3329) ;
                                                                                                                                           mul_add[1][50]<=((mult_out_10[50] + mult_out_11[50] + mult_out_12[50])%3329) ;
                                                                                                                                           mul_add[1][51]<=((mult_out_10[51] + mult_out_11[51] + mult_out_12[51])%3329) ;
                                                                                                                                           mul_add[1][52]<=((mult_out_10[52] + mult_out_11[52] + mult_out_12[52])%3329) ;
                                                                                                                                           mul_add[1][53]<=((mult_out_10[53] + mult_out_11[53] + mult_out_12[53])%3329) ;
                                                                                                                                           mul_add[1][54]<=((mult_out_10[54] + mult_out_11[54] + mult_out_12[54])%3329) ;
                                                                                                                                           mul_add[1][55]<=((mult_out_10[55] + mult_out_11[55] + mult_out_12[55])%3329) ;
                                                                                                                                           mul_add[1][56]<=((mult_out_10[56] + mult_out_11[56] + mult_out_12[56])%3329) ;
                                                                                                                                           mul_add[1][57]<=((mult_out_10[57] + mult_out_11[57] + mult_out_12[57])%3329) ;
                                                                                                                                           mul_add[1][58]<=((mult_out_10[58] + mult_out_11[58] + mult_out_12[58])%3329) ;
                                                                                                                                           mul_add[1][59]<=((mult_out_10[59] + mult_out_11[59] + mult_out_12[59])%3329) ;
                                                                                                                                           mul_add[1][60]<=((mult_out_10[60] + mult_out_11[60] + mult_out_12[60])%3329) ;
                                                                                                                                           mul_add[1][61]<=((mult_out_10[61] + mult_out_11[61] + mult_out_12[61])%3329) ;
                                                                                                                                           mul_add[1][62]<=((mult_out_10[62] + mult_out_11[62] + mult_out_12[62])%3329) ;
                                                                                                                                           mul_add[1][63]<=((mult_out_10[63] + mult_out_11[63] + mult_out_12[63])%3329) ;
                                                                                                                                           mul_add[1][64]<=((mult_out_10[64] + mult_out_11[64] + mult_out_12[64])%3329) ;
                                                                                                                                           mul_add[1][65]<=((mult_out_10[65] + mult_out_11[65] + mult_out_12[65])%3329) ;
                                                                                                                                           mul_add[1][66]<=((mult_out_10[66] + mult_out_11[66] + mult_out_12[66])%3329) ;
                                                                                                                                           mul_add[1][67]<=((mult_out_10[67] + mult_out_11[67] + mult_out_12[67])%3329) ;
                                                                                                                                           mul_add[1][68]<=((mult_out_10[68] + mult_out_11[68] + mult_out_12[68])%3329) ;
                                                                                                                                           mul_add[1][69]<=((mult_out_10[69] + mult_out_11[69] + mult_out_12[69])%3329) ;
                                                                                                                                           mul_add[1][70]<=((mult_out_10[70] + mult_out_11[70] + mult_out_12[70])%3329) ;
                                                                                                                                           mul_add[1][71]<=((mult_out_10[71] + mult_out_11[71] + mult_out_12[71])%3329) ;
                                                                                                                                           mul_add[1][72]<=((mult_out_10[72] + mult_out_11[72] + mult_out_12[72])%3329) ;
                                                                                                                                           mul_add[1][73]<=((mult_out_10[73] + mult_out_11[73] + mult_out_12[73])%3329) ;
                                                                                                                                           mul_add[1][74]<=((mult_out_10[74] + mult_out_11[74] + mult_out_12[74])%3329) ;
                                                                                                                                           mul_add[1][75]<=((mult_out_10[75] + mult_out_11[75] + mult_out_12[75])%3329) ;
                                                                                                                                           mul_add[1][76]<=((mult_out_10[76] + mult_out_11[76] + mult_out_12[76])%3329) ;
                                                                                                                                           mul_add[1][77]<=((mult_out_10[77] + mult_out_11[77] + mult_out_12[77])%3329) ;
                                                                                                                                           mul_add[1][78]<=((mult_out_10[78] + mult_out_11[78] + mult_out_12[78])%3329) ;
                                                                                                                                           mul_add[1][79]<=((mult_out_10[79] + mult_out_11[79] + mult_out_12[79])%3329) ;
                                                                                                                                           mul_add[1][80]<=((mult_out_10[80] + mult_out_11[80] + mult_out_12[80])%3329) ;
                                                                                                                                           mul_add[1][81]<=((mult_out_10[81] + mult_out_11[81] + mult_out_12[81])%3329) ;
                                                                                                                                           mul_add[1][82]<=((mult_out_10[82] + mult_out_11[82] + mult_out_12[82])%3329) ;
                                                                                                                                           mul_add[1][83]<=((mult_out_10[83] + mult_out_11[83] + mult_out_12[83])%3329) ;
                                                                                                                                           mul_add[1][84]<=((mult_out_10[84] + mult_out_11[84] + mult_out_12[84])%3329) ;
                                                                                                                                           mul_add[1][85]<=((mult_out_10[85] + mult_out_11[85] + mult_out_12[85])%3329) ;
                                                                                                                                           mul_add[1][86]<=((mult_out_10[86] + mult_out_11[86] + mult_out_12[86])%3329) ;
                                                                                                                                           mul_add[1][87]<=((mult_out_10[87] + mult_out_11[87] + mult_out_12[87])%3329) ;
                                                                                                                                           mul_add[1][88]<=((mult_out_10[88] + mult_out_11[88] + mult_out_12[88])%3329) ;
                                                                                                                                           mul_add[1][89]<=((mult_out_10[89] + mult_out_11[89] + mult_out_12[89])%3329) ;
                                                                                                                                           mul_add[1][90]<=((mult_out_10[90] + mult_out_11[90] + mult_out_12[90])%3329) ;
                                                                                                                                           mul_add[1][91]<=((mult_out_10[91] + mult_out_11[91] + mult_out_12[91])%3329) ;
                                                                                                                                           mul_add[1][92]<=((mult_out_10[92] + mult_out_11[92] + mult_out_12[92])%3329) ;
                                                                                                                                           mul_add[1][93]<=((mult_out_10[93] + mult_out_11[93] + mult_out_12[93])%3329) ;
                                                                                                                                           mul_add[1][94]<=((mult_out_10[94] + mult_out_11[94] + mult_out_12[94])%3329) ;
                                                                                                                                           mul_add[1][95]<=((mult_out_10[95] + mult_out_11[95] + mult_out_12[95])%3329) ;
                                                                                                                                           mul_add[1][96]<=((mult_out_10[96] + mult_out_11[96] + mult_out_12[96])%3329) ;
                                                                                                                                           mul_add[1][97]<=((mult_out_10[97] + mult_out_11[97] + mult_out_12[97])%3329) ;
                                                                                                                                           mul_add[1][98]<=((mult_out_10[98] + mult_out_11[98] + mult_out_12[98])%3329) ;
                                                                                                                                           mul_add[1][99]<=((mult_out_10[99] + mult_out_11[99] + mult_out_12[99])%3329) ;
                                                                                                                                           mul_add[1][100]<=((mult_out_10[100] + mult_out_11[100] + mult_out_12[100])%3329);
                                                                                                                                           mul_add[1][101]<=((mult_out_10[101] + mult_out_11[101] + mult_out_12[101])%3329) ;
                                                                                                                                           mul_add[1][102]<=((mult_out_10[102] + mult_out_11[102] + mult_out_12[102])%3329) ;
                                                                                                                                           mul_add[1][103]<=((mult_out_10[103] + mult_out_11[103] + mult_out_12[103])%3329) ;
                                                                                                                                           mul_add[1][104]<=((mult_out_10[104] + mult_out_11[104] + mult_out_12[104])%3329) ;
                                                                                                                                           mul_add[1][105]<=((mult_out_10[105] + mult_out_11[105] + mult_out_12[105])%3329) ;
                                                                                                                                           mul_add[1][106]<=((mult_out_10[106] + mult_out_11[106] + mult_out_12[106])%3329) ;
                                                                                                                                           mul_add[1][107]<=((mult_out_10[107] + mult_out_11[107] + mult_out_12[107])%3329) ;
                                                                                                                                           mul_add[1][108]<=((mult_out_10[108] + mult_out_11[108] + mult_out_12[108])%3329) ;
                                                                                                                                           mul_add[1][109]<=((mult_out_10[109] + mult_out_11[109] + mult_out_12[109])%3329) ;
                                                                                                                                           mul_add[1][110]<=((mult_out_10[110] + mult_out_11[110] + mult_out_12[110])%3329) ;
                                                                                                                                           mul_add[1][111]<=((mult_out_10[111] + mult_out_11[111] + mult_out_12[111])%3329) ;
                                                                                                                                           mul_add[1][112]<=((mult_out_10[112] + mult_out_11[112] + mult_out_12[112])%3329) ;
                                                                                                                                           mul_add[1][113]<=((mult_out_10[113] + mult_out_11[113] + mult_out_12[113])%3329) ;
                                                                                                                                           mul_add[1][114]<=((mult_out_10[114] + mult_out_11[114] + mult_out_12[114])%3329) ;
                                                                                                                                           mul_add[1][115]<=((mult_out_10[115] + mult_out_11[115] + mult_out_12[115])%3329) ;
                                                                                                                                           mul_add[1][116]<=((mult_out_10[116] + mult_out_11[116] + mult_out_12[116])%3329) ;
                                                                                                                                           mul_add[1][117]<=((mult_out_10[117] + mult_out_11[117] + mult_out_12[117])%3329) ;
                                                                                                                                           mul_add[1][118]<=((mult_out_10[118] + mult_out_11[118] + mult_out_12[118])%3329) ;
                                                                                                                                           mul_add[1][119]<=((mult_out_10[119] + mult_out_11[119] + mult_out_12[119])%3329) ;
                                                                                                                                           mul_add[1][120]<=((mult_out_10[120] + mult_out_11[120] + mult_out_12[120])%3329) ;
                                                                                                                                           mul_add[1][121]<=((mult_out_10[121] + mult_out_11[121] + mult_out_12[121])%3329) ;
                                                                                                                                           mul_add[1][122]<=((mult_out_10[122] + mult_out_11[122] + mult_out_12[122])%3329) ;
                                                                                                                                           mul_add[1][123]<=((mult_out_10[123] + mult_out_11[123] + mult_out_12[123])%3329);
                                                                                                                                           mul_add[1][124]<=((mult_out_10[124] + mult_out_11[124] + mult_out_12[124])%3329);
                                                                                                                                           mul_add[1][125]<=((mult_out_10[125] + mult_out_11[125] + mult_out_12[125])%3329);
                                                                                                                                           mul_add[1][126]<=((mult_out_10[126] + mult_out_11[126] + mult_out_12[126])%3329);
                                                                                                                                           mul_add[1][127]<=((mult_out_10[127] + mult_out_11[127] + mult_out_12[127])%3329);
                                                                                                                                           mul_add[1][128]<=((mult_out_10[128] + mult_out_11[128] + mult_out_12[128])%3329);
                                                                                                                                           mul_add[1][129]<=((mult_out_10[129] + mult_out_11[129] + mult_out_12[129])%3329);
                                                                                                                                           mul_add[1][130]<=((mult_out_10[130] + mult_out_11[130] + mult_out_12[130])%3329);
                                                                                                                                           mul_add[1][131]<=((mult_out_10[131] + mult_out_11[131] + mult_out_12[131])%3329);
                                                                                                                                           mul_add[1][132]<=((mult_out_10[132] + mult_out_11[132] + mult_out_12[132])%3329);
                                                                                                                                           mul_add[1][133]<=((mult_out_10[133] + mult_out_11[133] + mult_out_12[133])%3329);
                                                                                                                                           mul_add[1][134]<=((mult_out_10[134] + mult_out_11[134] + mult_out_12[134])%3329);
                                                                                                                                           mul_add[1][135]<=((mult_out_10[135] + mult_out_11[135] + mult_out_12[135])%3329);
                                                                                                                                           mul_add[1][136]<=((mult_out_10[136] + mult_out_11[136] + mult_out_12[136])%3329);
                                                                                                                                           mul_add[1][137]<=((mult_out_10[137] + mult_out_11[137] + mult_out_12[137])%3329);
                                                                                                                                           mul_add[1][138]<=((mult_out_10[138] + mult_out_11[138] + mult_out_12[138])%3329);
                                                                                                                                           mul_add[1][139]<=((mult_out_10[139] + mult_out_11[139] + mult_out_12[139])%3329);
                                                                                                                                           mul_add[1][140]<=((mult_out_10[140] + mult_out_11[140] + mult_out_12[140])%3329);
                                                                                                                                           mul_add[1][141]<=((mult_out_10[141] + mult_out_11[141] + mult_out_12[141])%3329);
                                                                                                                                           mul_add[1][142]<=((mult_out_10[142] + mult_out_11[142] + mult_out_12[142])%3329);
                                                                                                                                           mul_add[1][143]<=((mult_out_10[143] + mult_out_11[143] + mult_out_12[143])%3329);
                                                                                                                                           mul_add[1][144]<=((mult_out_10[144] + mult_out_11[144] + mult_out_12[144])%3329);
                                                                                                                                           mul_add[1][145]<=((mult_out_10[145] + mult_out_11[145] + mult_out_12[145])%3329);
                                                                                                                                           mul_add[1][146]<=((mult_out_10[146] + mult_out_11[146] + mult_out_12[146])%3329);
                                                                                                                                           mul_add[1][147]<=((mult_out_10[147] + mult_out_11[147] + mult_out_12[147])%3329);
                                                                                                                                           mul_add[1][148]<=((mult_out_10[148] + mult_out_11[148] + mult_out_12[148])%3329);
                                                                                                                                           mul_add[1][149]<=((mult_out_10[149] + mult_out_11[149] + mult_out_12[149])%3329);
                                                                                                                                           mul_add[1][150]<=((mult_out_10[150] + mult_out_11[150] + mult_out_12[150])%3329);
                                                                                                                                           mul_add[1][151]<=((mult_out_10[151] + mult_out_11[151] + mult_out_12[151])%3329);
                                                                                                                                           mul_add[1][152]<=((mult_out_10[152] + mult_out_11[152] + mult_out_12[152])%3329);
                                                                                                                                           mul_add[1][153]<=((mult_out_10[153] + mult_out_11[153] + mult_out_12[153])%3329);
                                                                                                                                           mul_add[1][154]<=((mult_out_10[154] + mult_out_11[154] + mult_out_12[154])%3329);
                                                                                                                                           mul_add[1][155]<=((mult_out_10[155] + mult_out_11[155] + mult_out_12[155])%3329);
                                                                                                                                           mul_add[1][156]<=((mult_out_10[156] + mult_out_11[156] + mult_out_12[156])%3329);
                                                                                                                                           mul_add[1][157]<=((mult_out_10[157] + mult_out_11[157] + mult_out_12[157])%3329) ;
                                                                                                                                           mul_add[1][158]<=((mult_out_10[158] + mult_out_11[158] + mult_out_12[158])%3329) ;
                                                                                                                                           mul_add[1][159]<=((mult_out_10[159] + mult_out_11[159] + mult_out_12[159])%3329);
                                                                                                                                           mul_add[1][160]<=((mult_out_10[160] + mult_out_11[160] + mult_out_12[160])%3329) ;
                                                                                                                                           mul_add[1][161]<=((mult_out_10[161] + mult_out_11[161] + mult_out_12[161])%3329) ;
                                                                                                                                           mul_add[1][162]<=((mult_out_10[162] + mult_out_11[162] + mult_out_12[162])%3329) ;
                                                                                                                                           mul_add[1][163]<=((mult_out_10[163] + mult_out_11[163] + mult_out_12[163])%3329);
                                                                                                                                           mul_add[1][164]<=((mult_out_10[164] + mult_out_11[164] + mult_out_12[164])%3329);
                                                                                                                                           mul_add[1][165]<=((mult_out_10[165] + mult_out_11[165] + mult_out_12[165])%3329) ;
                                                                                                                                           mul_add[1][166]<=((mult_out_10[166] + mult_out_11[166] + mult_out_12[166])%3329) ;
                                                                                                                                           mul_add[1][167]<=((mult_out_10[167] + mult_out_11[167] + mult_out_12[167])%3329) ;
                                                                                                                                           mul_add[1][168]<=((mult_out_10[168] + mult_out_11[168] + mult_out_12[168])%3329) ;
                                                                                                                                           mul_add[1][169]<=((mult_out_10[169] + mult_out_11[169] + mult_out_12[169])%3329) ;
                                                                                                                                           mul_add[1][170]<=((mult_out_10[170] + mult_out_11[170] + mult_out_12[170])%3329) ;
                                                                                                                                           mul_add[1][171]<=((mult_out_10[171] + mult_out_11[171] + mult_out_12[171])%3329) ;
                                                                                                                                           mul_add[1][172]<=((mult_out_10[172] + mult_out_11[172] + mult_out_12[172])%3329) ;
                                                                                                                                           mul_add[1][173]<=((mult_out_10[173] + mult_out_11[173] + mult_out_12[173])%3329) ;
                                                                                                                                           mul_add[1][174]<=((mult_out_10[174] + mult_out_11[174] + mult_out_12[174])%3329) ;
                                                                                                                                           mul_add[1][175]<=((mult_out_10[175] + mult_out_11[175] + mult_out_12[175])%3329) ;
                                                                                                                                           mul_add[1][176]<=((mult_out_10[176] + mult_out_11[176] + mult_out_12[176])%3329) ;
                                                                                                                                           mul_add[1][177]<=((mult_out_10[177] + mult_out_11[177] + mult_out_12[177])%3329) ;
                                                                                                                                           mul_add[1][178]<=((mult_out_10[178] + mult_out_11[178] + mult_out_12[178])%3329) ;
                                                                                                                                           mul_add[1][179]<=((mult_out_10[179] + mult_out_11[179] + mult_out_12[179])%3329) ;
                                                                                                                                           mul_add[1][180]<=((mult_out_10[180] + mult_out_11[180] + mult_out_12[180])%3329) ;
                                                                                                                                           mul_add[1][181]<=((mult_out_10[181] + mult_out_11[181] + mult_out_12[181])%3329) ;
                                                                                                                                           mul_add[1][182]<=((mult_out_10[182] + mult_out_11[182] + mult_out_12[182])%3329) ;
                                                                                                                                           mul_add[1][183]<=((mult_out_10[183] + mult_out_11[183] + mult_out_12[183])%3329) ;
                                                                                                                                           mul_add[1][184]<=((mult_out_10[184] + mult_out_11[184] + mult_out_12[184])%3329) ;
                                                                                                                                           mul_add[1][185]<=((mult_out_10[185] + mult_out_11[185] + mult_out_12[185])%3329) ;
                                                                                                                                           mul_add[1][186]<=((mult_out_10[186] + mult_out_11[186] + mult_out_12[186])%3329) ;
                                                                                                                                           mul_add[1][187]<=((mult_out_10[187] + mult_out_11[187] + mult_out_12[187])%3329) ;
                                                                                                                                           mul_add[1][188]<=((mult_out_10[188] + mult_out_11[188] + mult_out_12[188])%3329) ;
                                                                                                                                           mul_add[1][189]<=((mult_out_10[189] + mult_out_11[189] + mult_out_12[189])%3329) ;
                                                                                                                                           mul_add[1][190]<=((mult_out_10[190] + mult_out_11[190] + mult_out_12[190])%3329) ;
                                                                                                                                           mul_add[1][191]<=((mult_out_10[191] + mult_out_11[191] + mult_out_12[191])%3329) ;
                                                                                                                                           mul_add[1][192]<=((mult_out_10[192] + mult_out_11[192] + mult_out_12[192])%3329) ;
                                                                                                                                           mul_add[1][193]<=((mult_out_10[193] + mult_out_11[193] + mult_out_12[193])%3329) ;
                                                                                                                                           mul_add[1][194]<=((mult_out_10[194] + mult_out_11[194] + mult_out_12[194])%3329) ;
                                                                                                                                           mul_add[1][195]<=((mult_out_10[195] + mult_out_11[195] + mult_out_12[195])%3329) ;
                                                                                                                                           mul_add[1][196]<=((mult_out_10[196] + mult_out_11[196] + mult_out_12[196])%3329) ;
                                                                                                                                           mul_add[1][197]<=((mult_out_10[197] + mult_out_11[197] + mult_out_12[197])%3329) ;
                                                                                                                                           mul_add[1][198]<=((mult_out_10[198] + mult_out_11[198] + mult_out_12[198])%3329) ;
                                                                                                                                           mul_add[1][199]<=((mult_out_10[199] + mult_out_11[199] + mult_out_12[199])%3329) ;
                                                                                                                                           mul_add[1][200]<=((mult_out_10[200] + mult_out_11[200] + mult_out_12[200])%3329) ;
                                                                                                                                           mul_add[1][201]<=((mult_out_10[201] + mult_out_11[201] + mult_out_12[201])%3329) ;
                                                                                                                                           mul_add[1][202]<=((mult_out_10[202] + mult_out_11[202] + mult_out_12[202])%3329) ;
                                                                                                                                           mul_add[1][203]<=((mult_out_10[203] + mult_out_11[203] + mult_out_12[203])%3329) ;
                                                                                                                                           mul_add[1][204]<=((mult_out_10[204] + mult_out_11[204] + mult_out_12[204])%3329) ;
                                                                                                                                           mul_add[1][205]<=((mult_out_10[205] + mult_out_11[205] + mult_out_12[205])%3329) ;
                                                                                                                                           mul_add[1][206]<=((mult_out_10[206] + mult_out_11[206] + mult_out_12[206])%3329) ;
                                                                                                                                           mul_add[1][207]<=((mult_out_10[207] + mult_out_11[207] + mult_out_12[207])%3329) ;
                                                                                                                                           mul_add[1][208]<=((mult_out_10[208] + mult_out_11[208] + mult_out_12[208])%3329) ;
                                                                                                                                           mul_add[1][209]<=((mult_out_10[209] + mult_out_11[209] + mult_out_12[209])%3329) ;
                                                                                                                                           mul_add[1][210]<=((mult_out_10[210] + mult_out_11[210] + mult_out_12[210])%3329) ;
                                                                                                                                           mul_add[1][211]<=((mult_out_10[211] + mult_out_11[211] + mult_out_12[211])%3329) ;
                                                                                                                                           mul_add[1][212]<=((mult_out_10[212] + mult_out_11[212] + mult_out_12[212])%3329) ;
                                                                                                                                           mul_add[1][213]<=((mult_out_10[213] + mult_out_11[213] + mult_out_12[213])%3329) ;
                                                                                                                                           mul_add[1][214]<=((mult_out_10[214] + mult_out_11[214] + mult_out_12[214])%3329) ;
                                                                                                                                           mul_add[1][215]<=((mult_out_10[215] + mult_out_11[215] + mult_out_12[215])%3329) ;
                                                                                                                                           mul_add[1][216]<=((mult_out_10[216] + mult_out_11[216] + mult_out_12[216])%3329) ;
                                                                                                                                           mul_add[1][217]<=((mult_out_10[217] + mult_out_11[217] + mult_out_12[217])%3329) ;
                                                                                                                                           mul_add[1][218]<=((mult_out_10[218] + mult_out_11[218] + mult_out_12[218])%3329) ;
                                                                                                                                           mul_add[1][219]<=((mult_out_10[219] + mult_out_11[219] + mult_out_12[219])%3329) ;
                                                                                                                                           mul_add[1][220]<=((mult_out_10[220] + mult_out_11[220] + mult_out_12[220])%3329) ;
                                                                                                                                           mul_add[1][221]<=((mult_out_10[221] + mult_out_11[221] + mult_out_12[221])%3329) ;
                                                                                                                                           mul_add[1][222]<=((mult_out_10[222] + mult_out_11[222] + mult_out_12[222])%3329) ;
                                                                                                                                           mul_add[1][223]<=((mult_out_10[223] + mult_out_11[223] + mult_out_12[223])%3329) ;
                                                                                                                                           mul_add[1][224]<=((mult_out_10[224] + mult_out_11[224] + mult_out_12[224])%3329) ;
                                                                                                                                           mul_add[1][225]<=((mult_out_10[225] + mult_out_11[225] + mult_out_12[225])%3329) ;
                                                                                                                                           mul_add[1][226]<=((mult_out_10[226] + mult_out_11[226] + mult_out_12[226])%3329) ;
                                                                                                                                           mul_add[1][227]<=((mult_out_10[227] + mult_out_11[227] + mult_out_12[227])%3329) ;
                                                                                                                                           mul_add[1][228]<=((mult_out_10[228] + mult_out_11[228] + mult_out_12[228])%3329) ;
                                                                                                                                           mul_add[1][229]<=((mult_out_10[229] + mult_out_11[229] + mult_out_12[229])%3329) ;
                                                                                                                                           mul_add[1][230]<=((mult_out_10[230] + mult_out_11[230] + mult_out_12[230])%3329) ;
                                                                                                                                           mul_add[1][231]<=((mult_out_10[231] + mult_out_11[231] + mult_out_12[231])%3329) ;
                                                                                                                                           mul_add[1][232]<=((mult_out_10[232] + mult_out_11[232] + mult_out_12[232])%3329) ;
                                                                                                                                           mul_add[1][233]<=((mult_out_10[233] + mult_out_11[233] + mult_out_12[233])%3329) ;
                                                                                                                                           mul_add[1][234]<=((mult_out_10[234] + mult_out_11[234] + mult_out_12[234])%3329) ;
                                                                                                                                           mul_add[1][235]<=((mult_out_10[235] + mult_out_11[235] + mult_out_12[235])%3329) ;
                                                                                                                                           mul_add[1][236]<=((mult_out_10[236] + mult_out_11[236] + mult_out_12[236])%3329) ;
                                                                                                                                           mul_add[1][237]<=((mult_out_10[237] + mult_out_11[237] + mult_out_12[237])%3329) ;
                                                                                                                                           mul_add[1][238]<=((mult_out_10[238] + mult_out_11[238] + mult_out_12[238])%3329) ;
                                                                                                                                           mul_add[1][239]<=((mult_out_10[239] + mult_out_11[239] + mult_out_12[239])%3329) ;
                                                                                                                                           mul_add[1][240]<=((mult_out_10[240] + mult_out_11[240] + mult_out_12[240])%3329) ;
                                                                                                                                           mul_add[1][241]<=((mult_out_10[241] + mult_out_11[241] + mult_out_12[241])%3329) ;
                                                                                                                                           mul_add[1][242]<=((mult_out_10[242] + mult_out_11[242] + mult_out_12[242])%3329) ;
                                                                                                                                           mul_add[1][243]<=((mult_out_10[243] + mult_out_11[243] + mult_out_12[243])%3329) ;
                                                                                                                                           mul_add[1][244]<=((mult_out_10[244] + mult_out_11[244] + mult_out_12[244])%3329) ;
                                                                                                                                           mul_add[1][245]<=((mult_out_10[245] + mult_out_11[245] + mult_out_12[245])%3329) ;
                                                                                                                                           mul_add[1][246]<=((mult_out_10[246] + mult_out_11[246] + mult_out_12[246])%3329) ;
                                                                                                                                           mul_add[1][247]<=((mult_out_10[247] + mult_out_11[247] + mult_out_12[247])%3329);
                                                                                                                                           mul_add[1][248]<=((mult_out_10[248] + mult_out_11[248] + mult_out_12[248])%3329) ;
                                                                                                                                           mul_add[1][249]<=((mult_out_10[249] + mult_out_11[249] + mult_out_12[249])%3329) ;
                                                                                                                                           mul_add[1][250]<=((mult_out_10[250] + mult_out_11[250] + mult_out_12[250])%3329) ;
                                                                                                                                           mul_add[1][251]<=((mult_out_10[251] + mult_out_11[251] + mult_out_12[251])%3329) ;
                                                                                                                                           mul_add[1][252]<=((mult_out_10[252] + mult_out_11[252] + mult_out_12[252])%3329) ;
                                                                                                                                           mul_add[1][253]<=((mult_out_10[253] + mult_out_11[253] + mult_out_12[253])%3329) ;
                                                                                                                                           mul_add[1][254]<=((mult_out_10[254] + mult_out_11[254] + mult_out_12[254])%3329) ;
                                                                                                                                           mul_add[1][255]<=((mult_out_10[255] + mult_out_11[255] + mult_out_12[255])%3329) ;
                                                                                                                                          
                                                                                                                                      
                                                                                                                                           mul_add[2][0]<=((mult_out_20[0] + mult_out_21[0] + mult_out_22[0])%3329) ;
                                                                                                                                       mul_add[2][1]<=((mult_out_20[1] + mult_out_21[1] + mult_out_22[1])%3329) ;
                                                                                                                                       mul_add[2][2]<=((mult_out_20[2] + mult_out_21[2] + mult_out_22[2])%3329) ;
                                                                                                                                       mul_add[2][3]<=((mult_out_20[3] + mult_out_21[3] + mult_out_22[3])%3329) ;
                                                                                                                                       mul_add[2][4]<=((mult_out_20[4] + mult_out_21[4] + mult_out_22[4])%3329) ;
                                                                                                                                       mul_add[2][5]<=((mult_out_20[5] + mult_out_21[5] + mult_out_22[5])%3329) ;
                                                                                                                                       mul_add[2][6]<=((mult_out_20[6] + mult_out_21[6] + mult_out_22[6])%3329) ;
                                                                                                                                       mul_add[2][7]<=((mult_out_20[7] + mult_out_21[7] + mult_out_22[7])%3329) ;
                                                                                                                                       mul_add[2][8]<=((mult_out_20[8] + mult_out_21[8] + mult_out_22[8])%3329) ;
                                                                                                                                       mul_add[2][9]<=((mult_out_20[9] + mult_out_21[9] + mult_out_22[9])%3329) ;
                                                                                                                                       mul_add[2][10]<=((mult_out_20[10] + mult_out_21[10] + mult_out_22[10])%3329) ;
                                                                                                                                       mul_add[2][11]<=((mult_out_20[11] + mult_out_21[11] + mult_out_22[11])%3329) ;
                                                                                                                                       mul_add[2][12]<=((mult_out_20[12] + mult_out_21[12] + mult_out_22[12])%3329) ;
                                                                                                                                       mul_add[2][13]<=((mult_out_20[13] + mult_out_21[13] + mult_out_22[13])%3329) ;
                                                                                                                                       mul_add[2][14]<=((mult_out_20[14] + mult_out_21[14] + mult_out_22[14])%3329) ;
                                                                                                                                       mul_add[2][15]<=((mult_out_20[15] + mult_out_21[15] + mult_out_22[15])%3329) ;
                                                                                                                                       mul_add[2][16]<=((mult_out_20[16] + mult_out_21[16] + mult_out_22[16])%3329) ;
                                                                                                                                       mul_add[2][17]<=((mult_out_20[17] + mult_out_21[17] + mult_out_22[17])%3329) ;
                                                                                                                                       mul_add[2][18]<=((mult_out_20[18] + mult_out_21[18] + mult_out_22[18])%3329) ;
                                                                                                                                       mul_add[2][19]<=((mult_out_20[19] + mult_out_21[19] + mult_out_22[19])%3329) ;
                                                                                                                                       mul_add[2][20]<=((mult_out_20[20] + mult_out_21[20] + mult_out_22[20])%3329) ;
                                                                                                                                       mul_add[2][21]<=((mult_out_20[21] + mult_out_21[21] + mult_out_22[21])%3329) ;
                                                                                                                                       mul_add[2][22]<=((mult_out_20[22] + mult_out_21[22] + mult_out_22[22])%3329) ;
                                                                                                                                       mul_add[2][23]<=((mult_out_20[23] + mult_out_21[23] + mult_out_22[23])%3329) ;
                                                                                                                                       mul_add[2][24]<=((mult_out_20[24] + mult_out_21[24] + mult_out_22[24])%3329) ;
                                                                                                                                       mul_add[2][25]<=((mult_out_20[25] + mult_out_21[25] + mult_out_22[25])%3329) ;
                                                                                                                                       mul_add[2][26]<=((mult_out_20[26] + mult_out_21[26] + mult_out_22[26])%3329) ;
                                                                                                                                       mul_add[2][27]<=((mult_out_20[27] + mult_out_21[27] + mult_out_22[27])%3329) ;
                                                                                                                                       mul_add[2][28]<=((mult_out_20[28] + mult_out_21[28] + mult_out_22[28])%3329) ;
                                                                                                                                       mul_add[2][29]<=((mult_out_20[29] + mult_out_21[29] + mult_out_22[29])%3329) ;
                                                                                                                                       mul_add[2][30]<=((mult_out_20[30] + mult_out_21[30] + mult_out_22[30])%3329) ;
                                                                                                                                       mul_add[2][31]<=((mult_out_20[31] + mult_out_21[31] + mult_out_22[31])%3329) ;
                                                                                                                                       mul_add[2][32]<=((mult_out_20[32] + mult_out_21[32] + mult_out_22[32])%3329) ;
                                                                                                                                       mul_add[2][33]<=((mult_out_20[33] + mult_out_21[33] + mult_out_22[33])%3329) ;
                                                                                                                                       mul_add[2][34]<=((mult_out_20[34] + mult_out_21[34] + mult_out_22[34])%3329) ;
                                                                                                                                       mul_add[2][35]<=((mult_out_20[35] + mult_out_21[35] + mult_out_22[35])%3329) ;
                                                                                                                                       mul_add[2][36]<=((mult_out_20[36] + mult_out_21[36] + mult_out_22[36])%3329) ;
                                                                                                                                       mul_add[2][37]<=((mult_out_20[37] + mult_out_21[37] + mult_out_22[37])%3329) ;
                                                                                                                                       mul_add[2][38]<=((mult_out_20[38] + mult_out_21[38] + mult_out_22[38])%3329) ;
                                                                                                                                       mul_add[2][39]<=((mult_out_20[39] + mult_out_21[39] + mult_out_22[39])%3329) ;
                                                                                                                                       mul_add[2][40]<=((mult_out_20[40] + mult_out_21[40] + mult_out_22[40])%3329) ;
                                                                                                                                       mul_add[2][41]<=((mult_out_20[41] + mult_out_21[41] + mult_out_22[41])%3329) ;
                                                                                                                                       mul_add[2][42]<=((mult_out_20[42] + mult_out_21[42] + mult_out_22[42])%3329) ;
                                                                                                                                       mul_add[2][43]<=((mult_out_20[43] + mult_out_21[43] + mult_out_22[43])%3329) ;
                                                                                                                                       mul_add[2][44]<=((mult_out_20[44] + mult_out_21[44] + mult_out_22[44])%3329) ;
                                                                                                                                       mul_add[2][45]<=((mult_out_20[45] + mult_out_21[45] + mult_out_22[45])%3329) ;
                                                                                                                                       mul_add[2][46]<=((mult_out_20[46] + mult_out_21[46] + mult_out_22[46])%3329) ;
                                                                                                                                       mul_add[2][47]<=((mult_out_20[47] + mult_out_21[47] + mult_out_22[47])%3329) ;
                                                                                                                                       mul_add[2][48]<=((mult_out_20[48] + mult_out_21[48] + mult_out_22[48])%3329) ;
                                                                                                                                       mul_add[2][49]<=((mult_out_20[49] + mult_out_21[49] + mult_out_22[49])%3329) ;
                                                                                                                                       mul_add[2][50]<=((mult_out_20[50] + mult_out_21[50] + mult_out_22[50])%3329) ;
                                                                                                                                       mul_add[2][51]<=((mult_out_20[51] + mult_out_21[51] + mult_out_22[51])%3329) ;
                                                                                                                                       mul_add[2][52]<=((mult_out_20[52] + mult_out_21[52] + mult_out_22[52])%3329) ;
                                                                                                                                       mul_add[2][53]<=((mult_out_20[53] + mult_out_21[53] + mult_out_22[53])%3329) ;
                                                                                                                                       mul_add[2][54]<=((mult_out_20[54] + mult_out_21[54] + mult_out_22[54])%3329) ;
                                                                                                                                       mul_add[2][55]<=((mult_out_20[55] + mult_out_21[55] + mult_out_22[55])%3329) ;
                                                                                                                                       mul_add[2][56]<=((mult_out_20[56] + mult_out_21[56] + mult_out_22[56])%3329) ;
                                                                                                                                       mul_add[2][57]<=((mult_out_20[57] + mult_out_21[57] + mult_out_22[57])%3329) ;
                                                                                                                                       mul_add[2][58]<=((mult_out_20[58] + mult_out_21[58] + mult_out_22[58])%3329) ;
                                                                                                                                       mul_add[2][59]<=((mult_out_20[59] + mult_out_21[59] + mult_out_22[59])%3329) ;
                                                                                                                                       mul_add[2][60]<=((mult_out_20[60] + mult_out_21[60] + mult_out_22[60])%3329) ;
                                                                                                                                       mul_add[2][61]<=((mult_out_20[61] + mult_out_21[61] + mult_out_22[61])%3329) ;
                                                                                                                                       mul_add[2][62]<=((mult_out_20[62] + mult_out_21[62] + mult_out_22[62])%3329) ;
                                                                                                                                       mul_add[2][63]<=((mult_out_20[63] + mult_out_21[63] + mult_out_22[63])%3329) ;
                                                                                                                                       mul_add[2][64]<=((mult_out_20[64] + mult_out_21[64] + mult_out_22[64])%3329) ;
                                                                                                                                       mul_add[2][65]<=((mult_out_20[65] + mult_out_21[65] + mult_out_22[65])%3329) ;
                                                                                                                                       mul_add[2][66]<=((mult_out_20[66] + mult_out_21[66] + mult_out_22[66])%3329) ;
                                                                                                                                       mul_add[2][67]<=((mult_out_20[67] + mult_out_21[67] + mult_out_22[67])%3329) ;
                                                                                                                                       mul_add[2][68]<=((mult_out_20[68] + mult_out_21[68] + mult_out_22[68])%3329) ;
                                                                                                                                       mul_add[2][69]<=((mult_out_20[69] + mult_out_21[69] + mult_out_22[69])%3329) ;
                                                                                                                                       mul_add[2][70]<=((mult_out_20[70] + mult_out_21[70] + mult_out_22[70])%3329) ;
                                                                                                                                       mul_add[2][71]<=((mult_out_20[71] + mult_out_21[71] + mult_out_22[71])%3329) ;
                                                                                                                                       mul_add[2][72]<=((mult_out_20[72] + mult_out_21[72] + mult_out_22[72])%3329) ;
                                                                                                                                       mul_add[2][73]<=((mult_out_20[73] + mult_out_21[73] + mult_out_22[73])%3329) ;
                                                                                                                                       mul_add[2][74]<=((mult_out_20[74] + mult_out_21[74] + mult_out_22[74])%3329) ;
                                                                                                                                       mul_add[2][75]<=((mult_out_20[75] + mult_out_21[75] + mult_out_22[75])%3329) ;
                                                                                                                                       mul_add[2][76]<=((mult_out_20[76] + mult_out_21[76] + mult_out_22[76])%3329) ;
                                                                                                                                       mul_add[2][77]<=((mult_out_20[77] + mult_out_21[77] + mult_out_22[77])%3329) ;
                                                                                                                                       mul_add[2][78]<=((mult_out_20[78] + mult_out_21[78] + mult_out_22[78])%3329) ;
                                                                                                                                       mul_add[2][79]<=((mult_out_20[79] + mult_out_21[79] + mult_out_22[79])%3329) ;
                                                                                                                                       mul_add[2][80]<=((mult_out_20[80] + mult_out_21[80] + mult_out_22[80])%3329) ;
                                                                                                                                       mul_add[2][81]<=((mult_out_20[81] + mult_out_21[81] + mult_out_22[81])%3329) ;
                                                                                                                                       mul_add[2][82]<=((mult_out_20[82] + mult_out_21[82] + mult_out_22[82])%3329) ;
                                                                                                                                       mul_add[2][83]<=((mult_out_20[83] + mult_out_21[83] + mult_out_22[83])%3329) ;
                                                                                                                                       mul_add[2][84]<=((mult_out_20[84] + mult_out_21[84] + mult_out_22[84])%3329) ;
                                                                                                                                       mul_add[2][85]<=((mult_out_20[85] + mult_out_21[85] + mult_out_22[85])%3329) ;
                                                                                                                                       mul_add[2][86]<=((mult_out_20[86] + mult_out_21[86] + mult_out_22[86])%3329) ;
                                                                                                                                       mul_add[2][87]<=((mult_out_20[87] + mult_out_21[87] + mult_out_22[87])%3329) ;
                                                                                                                                       mul_add[2][88]<=((mult_out_20[88] + mult_out_21[88] + mult_out_22[88])%3329) ;
                                                                                                                                       mul_add[2][89]<=((mult_out_20[89] + mult_out_21[89] + mult_out_22[89])%3329) ;
                                                                                                                                       mul_add[2][90]<=((mult_out_20[90] + mult_out_21[90] + mult_out_22[90])%3329) ;
                                                                                                                                       mul_add[2][91]<=((mult_out_20[91] + mult_out_21[91] + mult_out_22[91])%3329) ;
                                                                                                                                       mul_add[2][92]<=((mult_out_20[92] + mult_out_21[92] + mult_out_22[92])%3329) ;
                                                                                                                                       mul_add[2][93]<=((mult_out_20[93] + mult_out_21[93] + mult_out_22[93])%3329) ;
                                                                                                                                       mul_add[2][94]<=((mult_out_20[94] + mult_out_21[94] + mult_out_22[94])%3329) ;
                                                                                                                                       mul_add[2][95]<=((mult_out_20[95] + mult_out_21[95] + mult_out_22[95])%3329) ;
                                                                                                                                       mul_add[2][96]<=((mult_out_20[96] + mult_out_21[96] + mult_out_22[96])%3329) ;
                                                                                                                                       mul_add[2][97]<=((mult_out_20[97] + mult_out_21[97] + mult_out_22[97])%3329) ;
                                                                                                                                       mul_add[2][98]<=((mult_out_20[98] + mult_out_21[98] + mult_out_22[98])%3329) ;
                                                                                                                                       mul_add[2][99]<=((mult_out_20[99] + mult_out_21[99] + mult_out_22[99])%3329) ;
                                                                                                                                       mul_add[2][100]<=((mult_out_20[100] + mult_out_21[100] + mult_out_22[100])%3329) ;
                                                                                                                                       mul_add[2][101]<=((mult_out_20[101] + mult_out_21[101] + mult_out_22[101])%3329) ;
                                                                                                                                       mul_add[2][102]<=((mult_out_20[102] + mult_out_21[102] + mult_out_22[102])%3329) ;
                                                                                                                                       mul_add[2][103]<=((mult_out_20[103] + mult_out_21[103] + mult_out_22[103])%3329) ;
                                                                                                                                       mul_add[2][104]<=((mult_out_20[104] + mult_out_21[104] + mult_out_22[104])%3329) ;
                                                                                                                                       mul_add[2][105]<=((mult_out_20[105] + mult_out_21[105] + mult_out_22[105])%3329) ;
                                                                                                                                       mul_add[2][106]<=((mult_out_20[106] + mult_out_21[106] + mult_out_22[106])%3329) ;
                                                                                                                                       mul_add[2][107]<=((mult_out_20[107] + mult_out_21[107] + mult_out_22[107])%3329) ;
                                                                                                                                       mul_add[2][108]<=((mult_out_20[108] + mult_out_21[108] + mult_out_22[108])%3329) ;
                                                                                                                                       mul_add[2][109]<=((mult_out_20[109] + mult_out_21[109] + mult_out_22[109])%3329) ;
                                                                                                                                       mul_add[2][110]<=((mult_out_20[110] + mult_out_21[110] + mult_out_22[110])%3329) ;
                                                                                                                                       mul_add[2][111]<=((mult_out_20[111] + mult_out_21[111] + mult_out_22[111])%3329) ;
                                                                                                                                       mul_add[2][112]<=((mult_out_20[112] + mult_out_21[112] + mult_out_22[112])%3329) ;
                                                                                                                                       mul_add[2][113]<=((mult_out_20[113] + mult_out_21[113] + mult_out_22[113])%3329) ;
                                                                                                                                       mul_add[2][114]<=((mult_out_20[114] + mult_out_21[114] + mult_out_22[114])%3329) ;
                                                                                                                                       mul_add[2][115]<=((mult_out_20[115] + mult_out_21[115] + mult_out_22[115])%3329) ;
                                                                                                                                       mul_add[2][116]<=((mult_out_20[116] + mult_out_21[116] + mult_out_22[116])%3329) ;
                                                                                                                                       mul_add[2][117]<=((mult_out_20[117] + mult_out_21[117] + mult_out_22[117])%3329) ;
                                                                                                                                       mul_add[2][118]<=((mult_out_20[118] + mult_out_21[118] + mult_out_22[118])%3329) ;
                                                                                                                                       mul_add[2][119]<=((mult_out_20[119] + mult_out_21[119] + mult_out_22[119])%3329) ;
                                                                                                                                       mul_add[2][120]<=((mult_out_20[120] + mult_out_21[120] + mult_out_22[120])%3329) ;
                                                                                                                                       mul_add[2][121]<=((mult_out_20[121] + mult_out_21[121] + mult_out_22[121])%3329) ;
                                                                                                                                       mul_add[2][122]<=((mult_out_20[122] + mult_out_21[122] + mult_out_22[122])%3329) ;
                                                                                                                                       mul_add[2][123]<=((mult_out_20[123] + mult_out_21[123] + mult_out_22[123])%3329) ;
                                                                                                                                       mul_add[2][124]<=((mult_out_20[124] + mult_out_21[124] + mult_out_22[124])%3329) ;
                                                                                                                                       mul_add[2][125]<=((mult_out_20[125] + mult_out_21[125] + mult_out_22[125])%3329) ;
                                                                                                                                       mul_add[2][126]<=((mult_out_20[126] + mult_out_21[126] + mult_out_22[126])%3329) ;
                                                                                                                                       mul_add[2][127]<=((mult_out_20[127] + mult_out_21[127] + mult_out_22[127])%3329) ;
                                                                                                                                       mul_add[2][128]<=((mult_out_20[128] + mult_out_21[128] + mult_out_22[128])%3329) ;
                                                                                                                                       mul_add[2][129]<=((mult_out_20[129] + mult_out_21[129] + mult_out_22[129])%3329) ;
                                                                                                                                       mul_add[2][130]<=((mult_out_20[130] + mult_out_21[130] + mult_out_22[130])%3329) ;
                                                                                                                                       mul_add[2][131]<=((mult_out_20[131] + mult_out_21[131] + mult_out_22[131])%3329) ;
                                                                                                                                       mul_add[2][132]<=((mult_out_20[132] + mult_out_21[132] + mult_out_22[132])%3329) ;
                                                                                                                                       mul_add[2][133]<=((mult_out_20[133] + mult_out_21[133] + mult_out_22[133])%3329) ;
                                                                                                                                       mul_add[2][134]<=((mult_out_20[134] + mult_out_21[134] + mult_out_22[134])%3329) ;
                                                                                                                                       mul_add[2][135]<=((mult_out_20[135] + mult_out_21[135] + mult_out_22[135])%3329) ;
                                                                                                                                       mul_add[2][136]<=((mult_out_20[136] + mult_out_21[136] + mult_out_22[136])%3329) ;
                                                                                                                                       mul_add[2][137]<=((mult_out_20[137] + mult_out_21[137] + mult_out_22[137])%3329) ;
                                                                                                                                       mul_add[2][138]<=((mult_out_20[138] + mult_out_21[138] + mult_out_22[138])%3329) ;
                                                                                                                                       mul_add[2][139]<=((mult_out_20[139] + mult_out_21[139] + mult_out_22[139])%3329) ;
                                                                                                                                       mul_add[2][140]<=((mult_out_20[140] + mult_out_21[140] + mult_out_22[140])%3329) ;
                                                                                                                                       mul_add[2][141]<=((mult_out_20[141] + mult_out_21[141] + mult_out_22[141])%3329) ;
                                                                                                                                       mul_add[2][142]<=((mult_out_20[142] + mult_out_21[142] + mult_out_22[142])%3329) ;
                                                                                                                                       mul_add[2][143]<=((mult_out_20[143] + mult_out_21[143] + mult_out_22[143])%3329) ;
                                                                                                                                       mul_add[2][144]<=((mult_out_20[144] + mult_out_21[144] + mult_out_22[144])%3329) ;
                                                                                                                                       mul_add[2][145]<=((mult_out_20[145] + mult_out_21[145] + mult_out_22[145])%3329) ;
                                                                                                                                       mul_add[2][146]<=((mult_out_20[146] + mult_out_21[146] + mult_out_22[146])%3329) ;
                                                                                                                                       mul_add[2][147]<=((mult_out_20[147] + mult_out_21[147] + mult_out_22[147])%3329) ;
                                                                                                                                       mul_add[2][148]<=((mult_out_20[148] + mult_out_21[148] + mult_out_22[148])%3329) ;
                                                                                                                                       mul_add[2][149]<=((mult_out_20[149] + mult_out_21[149] + mult_out_22[149])%3329) ;
                                                                                                                                       mul_add[2][150]<=((mult_out_20[150] + mult_out_21[150] + mult_out_22[150])%3329) ;
                                                                                                                                       mul_add[2][151]<=((mult_out_20[151] + mult_out_21[151] + mult_out_22[151])%3329) ;
                                                                                                                                       mul_add[2][152]<=((mult_out_20[152] + mult_out_21[152] + mult_out_22[152])%3329) ;
                                                                                                                                       mul_add[2][153]<=((mult_out_20[153] + mult_out_21[153] + mult_out_22[153])%3329) ;
                                                                                                                                       mul_add[2][154]<=((mult_out_20[154] + mult_out_21[154] + mult_out_22[154])%3329) ;
                                                                                                                                       mul_add[2][155]<=((mult_out_20[155] + mult_out_21[155] + mult_out_22[155])%3329) ;
                                                                                                                                       mul_add[2][156]<=((mult_out_20[156] + mult_out_21[156] + mult_out_22[156])%3329) ;
                                                                                                                                       mul_add[2][157]<=((mult_out_20[157] + mult_out_21[157] + mult_out_22[157])%3329) ;
                                                                                                                                       mul_add[2][158]<=((mult_out_20[158] + mult_out_21[158] + mult_out_22[158])%3329) ;
                                                                                                                                       mul_add[2][159]<=((mult_out_20[159] + mult_out_21[159] + mult_out_22[159])%3329) ;
                                                                                                                                       mul_add[2][160]<=((mult_out_20[160] + mult_out_21[160] + mult_out_22[160])%3329) ;
                                                                                                                                       mul_add[2][161]<=((mult_out_20[161] + mult_out_21[161] + mult_out_22[161])%3329) ;
                                                                                                                                       mul_add[2][162]<=((mult_out_20[162] + mult_out_21[162] + mult_out_22[162])%3329) ;
                                                                                                                                       mul_add[2][163]<=((mult_out_20[163] + mult_out_21[163] + mult_out_22[163])%3329) ;
                                                                                                                                       mul_add[2][164]<=((mult_out_20[164] + mult_out_21[164] + mult_out_22[164])%3329) ;
                                                                                                                                       mul_add[2][165]<=((mult_out_20[165] + mult_out_21[165] + mult_out_22[165])%3329) ;
                                                                                                                                       mul_add[2][166]<=((mult_out_20[166] + mult_out_21[166] + mult_out_22[166])%3329) ;
                                                                                                                                       mul_add[2][167]<=((mult_out_20[167] + mult_out_21[167] + mult_out_22[167])%3329) ;
                                                                                                                                       mul_add[2][168]<=((mult_out_20[168] + mult_out_21[168] + mult_out_22[168])%3329) ;
                                                                                                                                       mul_add[2][169]<=((mult_out_20[169] + mult_out_21[169] + mult_out_22[169])%3329) ;
                                                                                                                                       mul_add[2][170]<=((mult_out_20[170] + mult_out_21[170] + mult_out_22[170])%3329) ;
                                                                                                                                       mul_add[2][171]<=((mult_out_20[171] + mult_out_21[171] + mult_out_22[171])%3329) ;
                                                                                                                                       mul_add[2][172]<=((mult_out_20[172] + mult_out_21[172] + mult_out_22[172])%3329) ;
                                                                                                                                       mul_add[2][173]<=((mult_out_20[173] + mult_out_21[173] + mult_out_22[173])%3329) ;
                                                                                                                                       mul_add[2][174]<=((mult_out_20[174] + mult_out_21[174] + mult_out_22[174])%3329) ;
                                                                                                                                       mul_add[2][175]<=((mult_out_20[175] + mult_out_21[175] + mult_out_22[175])%3329) ;
                                                                                                                                       mul_add[2][176]<=((mult_out_20[176] + mult_out_21[176] + mult_out_22[176])%3329) ;
                                                                                                                                       mul_add[2][177]<=((mult_out_20[177] + mult_out_21[177] + mult_out_22[177])%3329) ;
                                                                                                                                       mul_add[2][178]<=((mult_out_20[178] + mult_out_21[178] + mult_out_22[178])%3329) ;
                                                                                                                                       mul_add[2][179]<=((mult_out_20[179] + mult_out_21[179] + mult_out_22[179])%3329) ;
                                                                                                                                       mul_add[2][180]<=((mult_out_20[180] + mult_out_21[180] + mult_out_22[180])%3329) ;
                                                                                                                                       mul_add[2][181]<=((mult_out_20[181] + mult_out_21[181] + mult_out_22[181])%3329) ;
                                                                                                                                       mul_add[2][182]<=((mult_out_20[182] + mult_out_21[182] + mult_out_22[182])%3329) ;
                                                                                                                                       mul_add[2][183]<=((mult_out_20[183] + mult_out_21[183] + mult_out_22[183])%3329) ;
                                                                                                                                       mul_add[2][184]<=((mult_out_20[184] + mult_out_21[184] + mult_out_22[184])%3329) ;
                                                                                                                                       mul_add[2][185]<=((mult_out_20[185] + mult_out_21[185] + mult_out_22[185])%3329) ;
                                                                                                                                       mul_add[2][186]<=((mult_out_20[186] + mult_out_21[186] + mult_out_22[186])%3329) ;
                                                                                                                                       mul_add[2][187]<=((mult_out_20[187] + mult_out_21[187] + mult_out_22[187])%3329) ;
                                                                                                                                       mul_add[2][188]<=((mult_out_20[188] + mult_out_21[188] + mult_out_22[188])%3329) ;
                                                                                                                                       mul_add[2][189]<=((mult_out_20[189] + mult_out_21[189] + mult_out_22[189])%3329) ;
                                                                                                                                       mul_add[2][190]<=((mult_out_20[190] + mult_out_21[190] + mult_out_22[190])%3329) ;
                                                                                                                                       mul_add[2][191]<=((mult_out_20[191] + mult_out_21[191] + mult_out_22[191])%3329) ;
                                                                                                                                       mul_add[2][192]<=((mult_out_20[192] + mult_out_21[192] + mult_out_22[192])%3329) ;
                                                                                                                                       mul_add[2][193]<=((mult_out_20[193] + mult_out_21[193] + mult_out_22[193])%3329) ;
                                                                                                                                       mul_add[2][194]<=((mult_out_20[194] + mult_out_21[194] + mult_out_22[194])%3329) ;
                                                                                                                                       mul_add[2][195]<=((mult_out_20[195] + mult_out_21[195] + mult_out_22[195])%3329) ;
                                                                                                                                       mul_add[2][196]<=((mult_out_20[196] + mult_out_21[196] + mult_out_22[196])%3329) ;
                                                                                                                                       mul_add[2][197]<=((mult_out_20[197] + mult_out_21[197] + mult_out_22[197])%3329) ;
                                                                                                                                       mul_add[2][198]<=((mult_out_20[198] + mult_out_21[198] + mult_out_22[198])%3329) ;
                                                                                                                                       mul_add[2][199]<=((mult_out_20[199] + mult_out_21[199] + mult_out_22[199])%3329) ;
                                                                                                                                       mul_add[2][200]<=((mult_out_20[200] + mult_out_21[200] + mult_out_22[200])%3329) ;
                                                                                                                                       mul_add[2][201]<=((mult_out_20[201] + mult_out_21[201] + mult_out_22[201])%3329) ;
                                                                                                                                       mul_add[2][202]<=((mult_out_20[202] + mult_out_21[202] + mult_out_22[202])%3329) ;
                                                                                                                                       mul_add[2][203]<=((mult_out_20[203] + mult_out_21[203] + mult_out_22[203])%3329) ;
                                                                                                                                       mul_add[2][204]<=((mult_out_20[204] + mult_out_21[204] + mult_out_22[204])%3329) ;
                                                                                                                                       mul_add[2][205]<=((mult_out_20[205] + mult_out_21[205] + mult_out_22[205])%3329) ;
                                                                                                                                       mul_add[2][206]<=((mult_out_20[206] + mult_out_21[206] + mult_out_22[206])%3329) ;
                                                                                                                                       mul_add[2][207]<=((mult_out_20[207] + mult_out_21[207] + mult_out_22[207])%3329) ;
                                                                                                                                       mul_add[2][208]<=((mult_out_20[208] + mult_out_21[208] + mult_out_22[208])%3329) ;
                                                                                                                                       mul_add[2][209]<=((mult_out_20[209] + mult_out_21[209] + mult_out_22[209])%3329) ;
                                                                                                                                       mul_add[2][210]<=((mult_out_20[210] + mult_out_21[210] + mult_out_22[210])%3329) ;
                                                                                                                                       mul_add[2][211]<=((mult_out_20[211] + mult_out_21[211] + mult_out_22[211])%3329) ;
                                                                                                                                       mul_add[2][212]<=((mult_out_20[212] + mult_out_21[212] + mult_out_22[212])%3329) ;
                                                                                                                                       mul_add[2][213]<=((mult_out_20[213] + mult_out_21[213] + mult_out_22[213])%3329) ;
                                                                                                                                       mul_add[2][214]<=((mult_out_20[214] + mult_out_21[214] + mult_out_22[214])%3329) ;
                                                                                                                                       mul_add[2][215]<=((mult_out_20[215] + mult_out_21[215] + mult_out_22[215])%3329) ;
                                                                                                                                       mul_add[2][216]<=((mult_out_20[216] + mult_out_21[216] + mult_out_22[216])%3329) ;
                                                                                                                                       mul_add[2][217]<=((mult_out_20[217] + mult_out_21[217] + mult_out_22[217])%3329) ;
                                                                                                                                       mul_add[2][218]<=((mult_out_20[218] + mult_out_21[218] + mult_out_22[218])%3329) ;
                                                                                                                                       mul_add[2][219]<=((mult_out_20[219] + mult_out_21[219] + mult_out_22[219])%3329) ;
                                                                                                                                       mul_add[2][220]<=((mult_out_20[220] + mult_out_21[220] + mult_out_22[220])%3329) ;
                                                                                                                                       mul_add[2][221]<=((mult_out_20[221] + mult_out_21[221] + mult_out_22[221])%3329) ;
                                                                                                                                       mul_add[2][222]<=((mult_out_20[222] + mult_out_21[222] + mult_out_22[222])%3329) ;
                                                                                                                                       mul_add[2][223]<=((mult_out_20[223] + mult_out_21[223] + mult_out_22[223])%3329) ;
                                                                                                                                       mul_add[2][224]<=((mult_out_20[224] + mult_out_21[224] + mult_out_22[224])%3329) ;
                                                                                                                                       mul_add[2][225]<=((mult_out_20[225] + mult_out_21[225] + mult_out_22[225])%3329) ;
                                                                                                                                       mul_add[2][226]<=((mult_out_20[226] + mult_out_21[226] + mult_out_22[226])%3329) ;
                                                                                                                                       mul_add[2][227]<=((mult_out_20[227] + mult_out_21[227] + mult_out_22[227])%3329) ;
                                                                                                                                       mul_add[2][228]<=((mult_out_20[228] + mult_out_21[228] + mult_out_22[228])%3329) ;
                                                                                                                                       mul_add[2][229]<=((mult_out_20[229] + mult_out_21[229] + mult_out_22[229])%3329) ;
                                                                                                                                       mul_add[2][230]<=((mult_out_20[230] + mult_out_21[230] + mult_out_22[230])%3329) ;
                                                                                                                                       mul_add[2][231]<=((mult_out_20[231] + mult_out_21[231] + mult_out_22[231])%3329) ;
                                                                                                                                       mul_add[2][232]<=((mult_out_20[232] + mult_out_21[232] + mult_out_22[232])%3329) ;
                                                                                                                                       mul_add[2][233]<=((mult_out_20[233] + mult_out_21[233] + mult_out_22[233])%3329) ;
                                                                                                                                       mul_add[2][234]<=((mult_out_20[234] + mult_out_21[234] + mult_out_22[234])%3329) ;
                                                                                                                                       mul_add[2][235]<=((mult_out_20[235] + mult_out_21[235] + mult_out_22[235])%3329) ;
                                                                                                                                       mul_add[2][236]<=((mult_out_20[236] + mult_out_21[236] + mult_out_22[236])%3329) ;
                                                                                                                                       mul_add[2][237]<=((mult_out_20[237] + mult_out_21[237] + mult_out_22[237])%3329) ;
                                                                                                                                       mul_add[2][238]<=((mult_out_20[238] + mult_out_21[238] + mult_out_22[238])%3329) ;
                                                                                                                                       mul_add[2][239]<=((mult_out_20[239] + mult_out_21[239] + mult_out_22[239])%3329) ;
                                                                                                                                       mul_add[2][240]<=((mult_out_20[240] + mult_out_21[240] + mult_out_22[240])%3329) ;
                                                                                                                                       mul_add[2][241]<=((mult_out_20[241] + mult_out_21[241] + mult_out_22[241])%3329) ;
                                                                                                                                       mul_add[2][242]<=((mult_out_20[242] + mult_out_21[242] + mult_out_22[242])%3329) ;
                                                                                                                                       mul_add[2][243]<=((mult_out_20[243] + mult_out_21[243] + mult_out_22[243])%3329) ;
                                                                                                                                       mul_add[2][244]<=((mult_out_20[244] + mult_out_21[244] + mult_out_22[244])%3329) ;
                                                                                                                                       mul_add[2][245]<=((mult_out_20[245] + mult_out_21[245] + mult_out_22[245])%3329) ;
                                                                                                                                       mul_add[2][246]<=((mult_out_20[246] + mult_out_21[246] + mult_out_22[246])%3329) ;
                                                                                                                                       mul_add[2][247]<=((mult_out_20[247] + mult_out_21[247] + mult_out_22[247])%3329) ;
                                                                                                                                       mul_add[2][248]<=((mult_out_20[248] + mult_out_21[248] + mult_out_22[248])%3329) ;
                                                                                                                                       mul_add[2][249]<=((mult_out_20[249] + mult_out_21[249] + mult_out_22[249])%3329) ;
                                                                                                                                       mul_add[2][250]<=((mult_out_20[250] + mult_out_21[250] + mult_out_22[250])%3329) ;
                                                                                                                                       mul_add[2][251]<=((mult_out_20[251] + mult_out_21[251] + mult_out_22[251])%3329) ;
                                                                                                                                       mul_add[2][252]<=((mult_out_20[252] + mult_out_21[252] + mult_out_22[252])%3329) ;
                                                                                                                                       mul_add[2][253]<=((mult_out_20[253] + mult_out_21[253] + mult_out_22[253])%3329) ;
                                                                                                                                       mul_add[2][254]<=((mult_out_20[254] + mult_out_21[254] + mult_out_22[254])%3329) ;
                                                                                                                                       mul_add[2][255]<=((mult_out_20[255] + mult_out_21[255] + mult_out_22[255])%3329) ;
                                                                                                                                                                                                             
                                                                                                                                                           if (done9_mul && done10_mul && done11_mul) begin
                                                                                                                                                                  mul_add_t[0][0] <= (mult_out_1[0] + mult_out_2[0] + mult_out_3[0]) % 3329;
                                                                                                                                                                  mul_add_t[0][1] <= (mult_out_1[1] + mult_out_2[1] + mult_out_3[1]) % 3329;
                                                                                                                                                                  mul_add_t[0][2] <= (mult_out_1[2] + mult_out_2[2] + mult_out_3[2]) % 3329;
                                                                                                                                                                  mul_add_t[0][3] <= (mult_out_1[3] + mult_out_2[3] + mult_out_3[3]) % 3329;
                                                                                                                                                                  mul_add_t[0][4] <= (mult_out_1[4] + mult_out_2[4] + mult_out_3[4]) % 3329;
                                                                                                                                                                  mul_add_t[0][5] <= (mult_out_1[5] + mult_out_2[5] + mult_out_3[5]) % 3329;
                                                                                                                                                                  mul_add_t[0][6] <= (mult_out_1[6] + mult_out_2[6] + mult_out_3[6]) % 3329;
                                                                                                                                                                  mul_add_t[0][7] <= (mult_out_1[7] + mult_out_2[7] + mult_out_3[7]) % 3329;
                                                                                                                                                                  mul_add_t[0][8] <= (mult_out_1[8] + mult_out_2[8] + mult_out_3[8]) % 3329;
                                                                                                                                                                  mul_add_t[0][9] <= (mult_out_1[9] + mult_out_2[9] + mult_out_3[9]) % 3329;
                                                                                                                                                                  mul_add_t[0][10] <= (mult_out_1[10] + mult_out_2[10] + mult_out_3[10]) % 3329;
                                                                                                                                                                  mul_add_t[0][11] <= (mult_out_1[11] + mult_out_2[11] + mult_out_3[11]) % 3329;
                                                                                                                                                                  mul_add_t[0][12] <= (mult_out_1[12] + mult_out_2[12] + mult_out_3[12]) % 3329;
                                                                                                                                                                  mul_add_t[0][13] <= (mult_out_1[13] + mult_out_2[13] + mult_out_3[13]) % 3329;
                                                                                                                                                                  mul_add_t[0][14] <= (mult_out_1[14] + mult_out_2[14] + mult_out_3[14]) % 3329;
                                                                                                                                                                  mul_add_t[0][15] <= (mult_out_1[15] + mult_out_2[15] + mult_out_3[15]) % 3329;
                                                                                                                                                                  mul_add_t[0][16] <= (mult_out_1[16] + mult_out_2[16] + mult_out_3[16]) % 3329;
                                                                                                                                                                  mul_add_t[0][17] <= (mult_out_1[17] + mult_out_2[17] + mult_out_3[17]) % 3329;
                                                                                                                                                                  mul_add_t[0][18] <= (mult_out_1[18] + mult_out_2[18] + mult_out_3[18]) % 3329;
                                                                                                                                                                  mul_add_t[0][19] <= (mult_out_1[19] + mult_out_2[19] + mult_out_3[19]) % 3329;
                                                                                                                                                                  mul_add_t[0][20] <= (mult_out_1[20] + mult_out_2[20] + mult_out_3[20]) % 3329;
                                                                                                                                                                  mul_add_t[0][21] <= (mult_out_1[21] + mult_out_2[21] + mult_out_3[21]) % 3329;
                                                                                                                                                                  mul_add_t[0][22] <= (mult_out_1[22] + mult_out_2[22] + mult_out_3[22]) % 3329;
                                                                                                                                                                  mul_add_t[0][23] <= (mult_out_1[23] + mult_out_2[23] + mult_out_3[23]) % 3329;
                                                                                                                                                                  mul_add_t[0][24] <= (mult_out_1[24] + mult_out_2[24] + mult_out_3[24]) % 3329;
                                                                                                                                                                  mul_add_t[0][25] <= (mult_out_1[25] + mult_out_2[25] + mult_out_3[25]) % 3329;
                                                                                                                                                                  mul_add_t[0][26] <= (mult_out_1[26] + mult_out_2[26] + mult_out_3[26]) % 3329;
                                                                                                                                                                  mul_add_t[0][27] <= (mult_out_1[27] + mult_out_2[27] + mult_out_3[27]) % 3329;
                                                                                                                                                                  mul_add_t[0][28] <= (mult_out_1[28] + mult_out_2[28] + mult_out_3[28]) % 3329;
                                                                                                                                                                  mul_add_t[0][29] <= (mult_out_1[29] + mult_out_2[29] + mult_out_3[29]) % 3329;
                                                                                                                                                                  mul_add_t[0][30] <= (mult_out_1[30] + mult_out_2[30] + mult_out_3[30]) % 3329;
                                                                                                                                                                  mul_add_t[0][31] <= (mult_out_1[31] + mult_out_2[31] + mult_out_3[31]) % 3329;
                                                                                                                                                                  mul_add_t[0][32] <= (mult_out_1[32] + mult_out_2[32] + mult_out_3[32]) % 3329;
                                                                                                                                                                  mul_add_t[0][33] <= (mult_out_1[33] + mult_out_2[33] + mult_out_3[33]) % 3329;
                                                                                                                                                                  mul_add_t[0][34] <= (mult_out_1[34] + mult_out_2[34] + mult_out_3[34]) % 3329;
                                                                                                                                                                  mul_add_t[0][35] <= (mult_out_1[35] + mult_out_2[35] + mult_out_3[35]) % 3329;
                                                                                                                                                                  mul_add_t[0][36] <= (mult_out_1[36] + mult_out_2[36] + mult_out_3[36]) % 3329;
                                                                                                                                                                  mul_add_t[0][37] <= (mult_out_1[37] + mult_out_2[37] + mult_out_3[37]) % 3329;
                                                                                                                                                                  mul_add_t[0][38] <= (mult_out_1[38] + mult_out_2[38] + mult_out_3[38]) % 3329;
                                                                                                                                                                  mul_add_t[0][39] <= (mult_out_1[39] + mult_out_2[39] + mult_out_3[39]) % 3329;
                                                                                                                                                                  mul_add_t[0][40] <= (mult_out_1[40] + mult_out_2[40] + mult_out_3[40]) % 3329;
                                                                                                                                                                  mul_add_t[0][41] <= (mult_out_1[41] + mult_out_2[41] + mult_out_3[41]) % 3329;
                                                                                                                                                                  mul_add_t[0][42] <= (mult_out_1[42] + mult_out_2[42] + mult_out_3[42]) % 3329;
                                                                                                                                                                  mul_add_t[0][43] <= (mult_out_1[43] + mult_out_2[43] + mult_out_3[43]) % 3329;
                                                                                                                                                                  mul_add_t[0][44] <= (mult_out_1[44] + mult_out_2[44] + mult_out_3[44]) % 3329;
                                                                                                                                                                  mul_add_t[0][45] <= (mult_out_1[45] + mult_out_2[45] + mult_out_3[45]) % 3329;
                                                                                                                                                                  mul_add_t[0][46] <= (mult_out_1[46] + mult_out_2[46] + mult_out_3[46]) % 3329;
                                                                                                                                                                  mul_add_t[0][47] <= (mult_out_1[47] + mult_out_2[47] + mult_out_3[47]) % 3329;
                                                                                                                                                                  mul_add_t[0][48] <= (mult_out_1[48] + mult_out_2[48] + mult_out_3[48]) % 3329;
                                                                                                                                                                  mul_add_t[0][49] <= (mult_out_1[49] + mult_out_2[49] + mult_out_3[49]) % 3329;
                                                                                                                                                                  mul_add_t[0][50] <= (mult_out_1[50] + mult_out_2[50] + mult_out_3[50]) % 3329;
                                                                                                                                                                  mul_add_t[0][51] <= (mult_out_1[51] + mult_out_2[51] + mult_out_3[51]) % 3329;
                                                                                                                                                                  mul_add_t[0][52] <= (mult_out_1[52] + mult_out_2[52] + mult_out_3[52]) % 3329;
                                                                                                                                                                  mul_add_t[0][53] <= (mult_out_1[53] + mult_out_2[53] + mult_out_3[53]) % 3329;
                                                                                                                                                                  mul_add_t[0][54] <= (mult_out_1[54] + mult_out_2[54] + mult_out_3[54]) % 3329;
                                                                                                                                                                  mul_add_t[0][55] <= (mult_out_1[55] + mult_out_2[55] + mult_out_3[55]) % 3329;
                                                                                                                                                                  mul_add_t[0][56] <= (mult_out_1[56] + mult_out_2[56] + mult_out_3[56]) % 3329;
                                                                                                                                                                  mul_add_t[0][57] <= (mult_out_1[57] + mult_out_2[57] + mult_out_3[57]) % 3329;
                                                                                                                                                                  mul_add_t[0][58] <= (mult_out_1[58] + mult_out_2[58] + mult_out_3[58]) % 3329;
                                                                                                                                                                  mul_add_t[0][59] <= (mult_out_1[59] + mult_out_2[59] + mult_out_3[59]) % 3329;
                                                                                                                                                                  mul_add_t[0][60] <= (mult_out_1[60] + mult_out_2[60] + mult_out_3[60]) % 3329;
                                                                                                                                                                  mul_add_t[0][61] <= (mult_out_1[61] + mult_out_2[61] + mult_out_3[61]) % 3329;
                                                                                                                                                                  mul_add_t[0][62] <= (mult_out_1[62] + mult_out_2[62] + mult_out_3[62]) % 3329;
                                                                                                                                                                  mul_add_t[0][63] <= (mult_out_1[63] + mult_out_2[63] + mult_out_3[63]) % 3329;
                                                                                                                                                                  mul_add_t[0][64] <= (mult_out_1[64] + mult_out_2[64] + mult_out_3[64]) % 3329;
                                                                                                                                                                  mul_add_t[0][65] <= (mult_out_1[65] + mult_out_2[65] + mult_out_3[65]) % 3329;
                                                                                                                                                                  mul_add_t[0][66] <= (mult_out_1[66] + mult_out_2[66] + mult_out_3[66]) % 3329;
                                                                                                                                                                  mul_add_t[0][67] <= (mult_out_1[67] + mult_out_2[67] + mult_out_3[67]) % 3329;
                                                                                                                                                                  mul_add_t[0][68] <= (mult_out_1[68] + mult_out_2[68] + mult_out_3[68]) % 3329;
                                                                                                                                                                  mul_add_t[0][69] <= (mult_out_1[69] + mult_out_2[69] + mult_out_3[69]) % 3329;
                                                                                                                                                                  mul_add_t[0][70] <= (mult_out_1[70] + mult_out_2[70] + mult_out_3[70]) % 3329;
                                                                                                                                                                  mul_add_t[0][71] <= (mult_out_1[71] + mult_out_2[71] + mult_out_3[71]) % 3329;
                                                                                                                                                                  mul_add_t[0][72] <= (mult_out_1[72] + mult_out_2[72] + mult_out_3[72]) % 3329;
                                                                                                                                                                  mul_add_t[0][73] <= (mult_out_1[73] + mult_out_2[73] + mult_out_3[73]) % 3329;
                                                                                                                                                                  mul_add_t[0][74] <= (mult_out_1[74] + mult_out_2[74] + mult_out_3[74]) % 3329;
                                                                                                                                                                  mul_add_t[0][75] <= (mult_out_1[75] + mult_out_2[75] + mult_out_3[75]) % 3329;
                                                                                                                                                                  mul_add_t[0][76] <= (mult_out_1[76] + mult_out_2[76] + mult_out_3[76]) % 3329;
                                                                                                                                                                  mul_add_t[0][77] <= (mult_out_1[77] + mult_out_2[77] + mult_out_3[77]) % 3329;
                                                                                                                                                                  mul_add_t[0][78] <= (mult_out_1[78] + mult_out_2[78] + mult_out_3[78]) % 3329;
                                                                                                                                                                  mul_add_t[0][79] <= (mult_out_1[79] + mult_out_2[79] + mult_out_3[79]) % 3329;
                                                                                                                                                                  mul_add_t[0][80] <= (mult_out_1[80] + mult_out_2[80] + mult_out_3[80]) % 3329;
                                                                                                                                                                  mul_add_t[0][81] <= (mult_out_1[81] + mult_out_2[81] + mult_out_3[81]) % 3329;
                                                                                                                                                                  mul_add_t[0][82] <= (mult_out_1[82] + mult_out_2[82] + mult_out_3[82]) % 3329;
                                                                                                                                                                  mul_add_t[0][83] <= (mult_out_1[83] + mult_out_2[83] + mult_out_3[83]) % 3329;
                                                                                                                                                                  mul_add_t[0][84] <= (mult_out_1[84] + mult_out_2[84] + mult_out_3[84]) % 3329;
                                                                                                                                                                  mul_add_t[0][85] <= (mult_out_1[85] + mult_out_2[85] + mult_out_3[85]) % 3329;
                                                                                                                                                                  mul_add_t[0][86] <= (mult_out_1[86] + mult_out_2[86] + mult_out_3[86]) % 3329;
                                                                                                                                                                  mul_add_t[0][87] <= (mult_out_1[87] + mult_out_2[87] + mult_out_3[87]) % 3329;
                                                                                                                                                                  mul_add_t[0][88] <= (mult_out_1[88] + mult_out_2[88] + mult_out_3[88]) % 3329;
                                                                                                                                                                  mul_add_t[0][89] <= (mult_out_1[89] + mult_out_2[89] + mult_out_3[89]) % 3329;
                                                                                                                                                                  mul_add_t[0][90] <= (mult_out_1[90] + mult_out_2[90] + mult_out_3[90]) % 3329;
                                                                                                                                                                  mul_add_t[0][91] <= (mult_out_1[91] + mult_out_2[91] + mult_out_3[91]) % 3329;
                                                                                                                                                                  mul_add_t[0][92] <= (mult_out_1[92] + mult_out_2[92] + mult_out_3[92]) % 3329;
                                                                                                                                                                  mul_add_t[0][93] <= (mult_out_1[93] + mult_out_2[93] + mult_out_3[93]) % 3329;
                                                                                                                                                                  mul_add_t[0][94] <= (mult_out_1[94] + mult_out_2[94] + mult_out_3[94]) % 3329;
                                                                                                                                                                  mul_add_t[0][95] <= (mult_out_1[95] + mult_out_2[95] + mult_out_3[95]) % 3329;
                                                                                                                                                                  mul_add_t[0][96] <= (mult_out_1[96] + mult_out_2[96] + mult_out_3[96]) % 3329;
                                                                                                                                                                  mul_add_t[0][97] <= (mult_out_1[97] + mult_out_2[97] + mult_out_3[97]) % 3329;
                                                                                                                                                                  mul_add_t[0][98] <= (mult_out_1[98] + mult_out_2[98] + mult_out_3[98]) % 3329;
                                                                                                                                                                  mul_add_t[0][99] <= (mult_out_1[99] + mult_out_2[99] + mult_out_3[99]) % 3329;
                                                                                                                                                                  mul_add_t[0][100] <= (mult_out_1[100] + mult_out_2[100] + mult_out_3[100]) % 3329;
                                                                                                                                                                  mul_add_t[0][101] <= (mult_out_1[101] + mult_out_2[101] + mult_out_3[101]) % 3329;
                                                                                                                                                                  mul_add_t[0][102] <= (mult_out_1[102] + mult_out_2[102] + mult_out_3[102]) % 3329;
                                                                                                                                                                  mul_add_t[0][103] <= (mult_out_1[103] + mult_out_2[103] + mult_out_3[103]) % 3329;
                                                                                                                                                                  mul_add_t[0][104] <= (mult_out_1[104] + mult_out_2[104] + mult_out_3[104]) % 3329;
                                                                                                                                                                  mul_add_t[0][105] <= (mult_out_1[105] + mult_out_2[105] + mult_out_3[105]) % 3329;
                                                                                                                                                                  mul_add_t[0][106] <= (mult_out_1[106] + mult_out_2[106] + mult_out_3[106]) % 3329;
                                                                                                                                                                  mul_add_t[0][107] <= (mult_out_1[107] + mult_out_2[107] + mult_out_3[107]) % 3329;
                                                                                                                                                                  mul_add_t[0][108] <= (mult_out_1[108] + mult_out_2[108] + mult_out_3[108]) % 3329;
                                                                                                                                                                  mul_add_t[0][109] <= (mult_out_1[109] + mult_out_2[109] + mult_out_3[109]) % 3329;
                                                                                                                                                                  mul_add_t[0][110] <= (mult_out_1[110] + mult_out_2[110] + mult_out_3[110]) % 3329;
                                                                                                                                                                  mul_add_t[0][111] <= (mult_out_1[111] + mult_out_2[111] + mult_out_3[111]) % 3329;
                                                                                                                                                                  mul_add_t[0][112] <= (mult_out_1[112] + mult_out_2[112] + mult_out_3[112]) % 3329;
                                                                                                                                                                  mul_add_t[0][113] <= (mult_out_1[113] + mult_out_2[113] + mult_out_3[113]) % 3329;
                                                                                                                                                                  mul_add_t[0][114] <= (mult_out_1[114] + mult_out_2[114] + mult_out_3[114]) % 3329;
                                                                                                                                                                  mul_add_t[0][115] <= (mult_out_1[115] + mult_out_2[115] + mult_out_3[115]) % 3329;
                                                                                                                                                                  mul_add_t[0][116] <= (mult_out_1[116] + mult_out_2[116] + mult_out_3[116]) % 3329;
                                                                                                                                                                  mul_add_t[0][117] <= (mult_out_1[117] + mult_out_2[117] + mult_out_3[117]) % 3329;
                                                                                                                                                                  mul_add_t[0][118] <= (mult_out_1[118] + mult_out_2[118] + mult_out_3[118]) % 3329;
                                                                                                                                                                  mul_add_t[0][119] <= (mult_out_1[119] + mult_out_2[119] + mult_out_3[119]) % 3329;
                                                                                                                                                                  mul_add_t[0][120] <= (mult_out_1[120] + mult_out_2[120] + mult_out_3[120]) % 3329;
                                                                                                                                                                  mul_add_t[0][121] <= (mult_out_1[121] + mult_out_2[121] + mult_out_3[121]) % 3329;
                                                                                                                                                                  mul_add_t[0][122] <= (mult_out_1[122] + mult_out_2[122] + mult_out_3[122]) % 3329;
                                                                                                                                                                  mul_add_t[0][123] <= (mult_out_1[123] + mult_out_2[123] + mult_out_3[123]) % 3329;
                                                                                                                                                                  mul_add_t[0][124] <= (mult_out_1[124] + mult_out_2[124] + mult_out_3[124]) % 3329;
                                                                                                                                                                  mul_add_t[0][125] <= (mult_out_1[125] + mult_out_2[125] + mult_out_3[125]) % 3329;
                                                                                                                                                                  mul_add_t[0][126] <= (mult_out_1[126] + mult_out_2[126] + mult_out_3[126]) % 3329;
                                                                                                                                                                  mul_add_t[0][127] <= (mult_out_1[127] + mult_out_2[127] + mult_out_3[127]) % 3329;
                                                                                                                                                                  mul_add_t[0][128] <= (mult_out_1[128] + mult_out_2[128] + mult_out_3[128]) % 3329;
                                                                                                                                                                  mul_add_t[0][129] <= (mult_out_1[129] + mult_out_2[129] + mult_out_3[129]) % 3329;
                                                                                                                                                                  mul_add_t[0][130] <= (mult_out_1[130] + mult_out_2[130] + mult_out_3[130]) % 3329;
                                                                                                                                                                  mul_add_t[0][131] <= (mult_out_1[131] + mult_out_2[131] + mult_out_3[131]) % 3329;
                                                                                                                                                                  mul_add_t[0][132] <= (mult_out_1[132] + mult_out_2[132] + mult_out_3[132]) % 3329;
                                                                                                                                                                  mul_add_t[0][133] <= (mult_out_1[133] + mult_out_2[133] + mult_out_3[133]) % 3329;
                                                                                                                                                                  mul_add_t[0][134] <= (mult_out_1[134] + mult_out_2[134] + mult_out_3[134]) % 3329;
                                                                                                                                                                  mul_add_t[0][135] <= (mult_out_1[135] + mult_out_2[135] + mult_out_3[135]) % 3329;
                                                                                                                                                                  mul_add_t[0][136] <= (mult_out_1[136] + mult_out_2[136] + mult_out_3[136]) % 3329;
                                                                                                                                                                  mul_add_t[0][137] <= (mult_out_1[137] + mult_out_2[137] + mult_out_3[137]) % 3329;
                                                                                                                                                                  mul_add_t[0][138] <= (mult_out_1[138] + mult_out_2[138] + mult_out_3[138]) % 3329;
                                                                                                                                                                  mul_add_t[0][139] <= (mult_out_1[139] + mult_out_2[139] + mult_out_3[139]) % 3329;
                                                                                                                                                                  mul_add_t[0][140] <= (mult_out_1[140] + mult_out_2[140] + mult_out_3[140]) % 3329;
                                                                                                                                                                  mul_add_t[0][141] <= (mult_out_1[141] + mult_out_2[141] + mult_out_3[141]) % 3329;
                                                                                                                                                                  mul_add_t[0][142] <= (mult_out_1[142] + mult_out_2[142] + mult_out_3[142]) % 3329;
                                                                                                                                                                  mul_add_t[0][143] <= (mult_out_1[143] + mult_out_2[143] + mult_out_3[143]) % 3329;
                                                                                                                                                                  mul_add_t[0][144] <= (mult_out_1[144] + mult_out_2[144] + mult_out_3[144]) % 3329;
                                                                                                                                                                  mul_add_t[0][145] <= (mult_out_1[145] + mult_out_2[145] + mult_out_3[145]) % 3329;
                                                                                                                                                                  mul_add_t[0][146] <= (mult_out_1[146] + mult_out_2[146] + mult_out_3[146]) % 3329;
                                                                                                                                                                  mul_add_t[0][147] <= (mult_out_1[147] + mult_out_2[147] + mult_out_3[147]) % 3329;
                                                                                                                                                                  mul_add_t[0][148] <= (mult_out_1[148] + mult_out_2[148] + mult_out_3[148]) % 3329;
                                                                                                                                                                  mul_add_t[0][149] <= (mult_out_1[149] + mult_out_2[149] + mult_out_3[149]) % 3329;
                                                                                                                                                                  mul_add_t[0][150] <= (mult_out_1[150] + mult_out_2[150] + mult_out_3[150]) % 3329;
                                                                                                                                                                  mul_add_t[0][151] <= (mult_out_1[151] + mult_out_2[151] + mult_out_3[151]) % 3329;
                                                                                                                                                                  mul_add_t[0][152] <= (mult_out_1[152] + mult_out_2[152] + mult_out_3[152]) % 3329;
                                                                                                                                                                  mul_add_t[0][153] <= (mult_out_1[153] + mult_out_2[153] + mult_out_3[153]) % 3329;
                                                                                                                                                                  mul_add_t[0][154] <= (mult_out_1[154] + mult_out_2[154] + mult_out_3[154]) % 3329;
                                                                                                                                                                  mul_add_t[0][155] <= (mult_out_1[155] + mult_out_2[155] + mult_out_3[155]) % 3329;
                                                                                                                                                                  mul_add_t[0][156] <= (mult_out_1[156] + mult_out_2[156] + mult_out_3[156]) % 3329;
                                                                                                                                                                  mul_add_t[0][157] <= (mult_out_1[157] + mult_out_2[157] + mult_out_3[157]) % 3329;
                                                                                                                                                                  mul_add_t[0][158] <= (mult_out_1[158] + mult_out_2[158] + mult_out_3[158]) % 3329;
                                                                                                                                                                  mul_add_t[0][159] <= (mult_out_1[159] + mult_out_2[159] + mult_out_3[159]) % 3329;
                                                                                                                                                                  mul_add_t[0][160] <= (mult_out_1[160] + mult_out_2[160] + mult_out_3[160]) % 3329;
                                                                                                                                                                  mul_add_t[0][161] <= (mult_out_1[161] + mult_out_2[161] + mult_out_3[161]) % 3329;
                                                                                                                                                                  mul_add_t[0][162] <= (mult_out_1[162] + mult_out_2[162] + mult_out_3[162]) % 3329;
                                                                                                                                                                  mul_add_t[0][163] <= (mult_out_1[163] + mult_out_2[163] + mult_out_3[163]) % 3329;
                                                                                                                                                                  mul_add_t[0][164] <= (mult_out_1[164] + mult_out_2[164] + mult_out_3[164]) % 3329;
                                                                                                                                                                  mul_add_t[0][165] <= (mult_out_1[165] + mult_out_2[165] + mult_out_3[165]) % 3329;
                                                                                                                                                                  mul_add_t[0][166] <= (mult_out_1[166] + mult_out_2[166] + mult_out_3[166]) % 3329;
                                                                                                                                                                  mul_add_t[0][167] <= (mult_out_1[167] + mult_out_2[167] + mult_out_3[167]) % 3329;
                                                                                                                                                                  mul_add_t[0][168] <= (mult_out_1[168] + mult_out_2[168] + mult_out_3[168]) % 3329;
                                                                                                                                                                  mul_add_t[0][169] <= (mult_out_1[169] + mult_out_2[169] + mult_out_3[169]) % 3329;
                                                                                                                                                                  mul_add_t[0][170] <= (mult_out_1[170] + mult_out_2[170] + mult_out_3[170]) % 3329;
                                                                                                                                                                  mul_add_t[0][171] <= (mult_out_1[171] + mult_out_2[171] + mult_out_3[171]) % 3329;
                                                                                                                                                                  mul_add_t[0][172] <= (mult_out_1[172] + mult_out_2[172] + mult_out_3[172]) % 3329;
                                                                                                                                                                  mul_add_t[0][173] <= (mult_out_1[173] + mult_out_2[173] + mult_out_3[173]) % 3329;
                                                                                                                                                                  mul_add_t[0][174] <= (mult_out_1[174] + mult_out_2[174] + mult_out_3[174]) % 3329;
                                                                                                                                                                  mul_add_t[0][175] <= (mult_out_1[175] + mult_out_2[175] + mult_out_3[175]) % 3329;
                                                                                                                                                                  mul_add_t[0][176] <= (mult_out_1[176] + mult_out_2[176] + mult_out_3[176]) % 3329;
                                                                                                                                                                  mul_add_t[0][177] <= (mult_out_1[177] + mult_out_2[177] + mult_out_3[177]) % 3329;
                                                                                                                                                                  mul_add_t[0][178] <= (mult_out_1[178] + mult_out_2[178] + mult_out_3[178]) % 3329;
                                                                                                                                                                  mul_add_t[0][179] <= (mult_out_1[179] + mult_out_2[179] + mult_out_3[179]) % 3329;
                                                                                                                                                                  mul_add_t[0][180] <= (mult_out_1[180] + mult_out_2[180] + mult_out_3[180]) % 3329;
                                                                                                                                                                  mul_add_t[0][181] <= (mult_out_1[181] + mult_out_2[181] + mult_out_3[181]) % 3329;
                                                                                                                                                                  mul_add_t[0][182] <= (mult_out_1[182] + mult_out_2[182] + mult_out_3[182]) % 3329;
                                                                                                                                                                  mul_add_t[0][183] <= (mult_out_1[183] + mult_out_2[183] + mult_out_3[183]) % 3329;
                                                                                                                                                                  mul_add_t[0][184] <= (mult_out_1[184] + mult_out_2[184] + mult_out_3[184]) % 3329;
                                                                                                                                                                  mul_add_t[0][185] <= (mult_out_1[185] + mult_out_2[185] + mult_out_3[185]) % 3329;
                                                                                                                                                                  mul_add_t[0][186] <= (mult_out_1[186] + mult_out_2[186] + mult_out_3[186]) % 3329;
                                                                                                                                                                  mul_add_t[0][187] <= (mult_out_1[187] + mult_out_2[187] + mult_out_3[187]) % 3329;
                                                                                                                                                                  mul_add_t[0][188] <= (mult_out_1[188] + mult_out_2[188] + mult_out_3[188]) % 3329;
                                                                                                                                                                  mul_add_t[0][189] <= (mult_out_1[189] + mult_out_2[189] + mult_out_3[189]) % 3329;
                                                                                                                                                                  mul_add_t[0][190] <= (mult_out_1[190] + mult_out_2[190] + mult_out_3[190]) % 3329;
                                                                                                                                                                  mul_add_t[0][191] <= (mult_out_1[191] + mult_out_2[191] + mult_out_3[191]) % 3329;
                                                                                                                                                                  mul_add_t[0][192] <= (mult_out_1[192] + mult_out_2[192] + mult_out_3[192]) % 3329;
                                                                                                                                                                  mul_add_t[0][193] <= (mult_out_1[193] + mult_out_2[193] + mult_out_3[193]) % 3329;
                                                                                                                                                                  mul_add_t[0][194] <= (mult_out_1[194] + mult_out_2[194] + mult_out_3[194]) % 3329;
                                                                                                                                                                  mul_add_t[0][195] <= (mult_out_1[195] + mult_out_2[195] + mult_out_3[195]) % 3329;
                                                                                                                                                                  mul_add_t[0][196] <= (mult_out_1[196] + mult_out_2[196] + mult_out_3[196]) % 3329;
                                                                                                                                                                  mul_add_t[0][197] <= (mult_out_1[197] + mult_out_2[197] + mult_out_3[197]) % 3329;
                                                                                                                                                                  mul_add_t[0][198] <= (mult_out_1[198] + mult_out_2[198] + mult_out_3[198]) % 3329;
                                                                                                                                                                  mul_add_t[0][199] <= (mult_out_1[199] + mult_out_2[199] + mult_out_3[199]) % 3329;
                                                                                                                                                                  mul_add_t[0][200] <= (mult_out_1[200] + mult_out_2[200] + mult_out_3[200]) % 3329;
                                                                                                                                                                  mul_add_t[0][201] <= (mult_out_1[201] + mult_out_2[201] + mult_out_3[201]) % 3329;
                                                                                                                                                                  mul_add_t[0][202] <= (mult_out_1[202] + mult_out_2[202] + mult_out_3[202]) % 3329;
                                                                                                                                                                  mul_add_t[0][203] <= (mult_out_1[203] + mult_out_2[203] + mult_out_3[203]) % 3329;
                                                                                                                                                                  mul_add_t[0][204] <= (mult_out_1[204] + mult_out_2[204] + mult_out_3[204]) % 3329;
                                                                                                                                                                  mul_add_t[0][205] <= (mult_out_1[205] + mult_out_2[205] + mult_out_3[205]) % 3329;
                                                                                                                                                                  mul_add_t[0][206] <= (mult_out_1[206] + mult_out_2[206] + mult_out_3[206]) % 3329;
                                                                                                                                                                  mul_add_t[0][207] <= (mult_out_1[207] + mult_out_2[207] + mult_out_3[207]) % 3329;
                                                                                                                                                                  mul_add_t[0][208] <= (mult_out_1[208] + mult_out_2[208] + mult_out_3[208]) % 3329;
                                                                                                                                                                  mul_add_t[0][209] <= (mult_out_1[209] + mult_out_2[209] + mult_out_3[209]) % 3329;
                                                                                                                                                                  mul_add_t[0][210] <= (mult_out_1[210] + mult_out_2[210] + mult_out_3[210]) % 3329;
                                                                                                                                                                  mul_add_t[0][211] <= (mult_out_1[211] + mult_out_2[211] + mult_out_3[211]) % 3329;
                                                                                                                                                                  mul_add_t[0][212] <= (mult_out_1[212] + mult_out_2[212] + mult_out_3[212]) % 3329;
                                                                                                                                                                  mul_add_t[0][213] <= (mult_out_1[213] + mult_out_2[213] + mult_out_3[213]) % 3329;
                                                                                                                                                                  mul_add_t[0][214] <= (mult_out_1[214] + mult_out_2[214] + mult_out_3[214]) % 3329;
                                                                                                                                                                  mul_add_t[0][215] <= (mult_out_1[215] + mult_out_2[215] + mult_out_3[215]) % 3329;
                                                                                                                                                                  mul_add_t[0][216] <= (mult_out_1[216] + mult_out_2[216] + mult_out_3[216]) % 3329;
                                                                                                                                                                  mul_add_t[0][217] <= (mult_out_1[217] + mult_out_2[217] + mult_out_3[217]) % 3329;
                                                                                                                                                                  mul_add_t[0][218] <= (mult_out_1[218] + mult_out_2[218] + mult_out_3[218]) % 3329;
                                                                                                                                                                  mul_add_t[0][219] <= (mult_out_1[219] + mult_out_2[219] + mult_out_3[219]) % 3329;
                                                                                                                                                                  mul_add_t[0][220] <= (mult_out_1[220] + mult_out_2[220] + mult_out_3[220]) % 3329;
                                                                                                                                                                  mul_add_t[0][221] <= (mult_out_1[221] + mult_out_2[221] + mult_out_3[221]) % 3329;
                                                                                                                                                                  mul_add_t[0][222] <= (mult_out_1[222] + mult_out_2[222] + mult_out_3[222]) % 3329;
                                                                                                                                                                  mul_add_t[0][223] <= (mult_out_1[223] + mult_out_2[223] + mult_out_3[223]) % 3329;
                                                                                                                                                                  mul_add_t[0][224] <= (mult_out_1[224] + mult_out_2[224] + mult_out_3[224]) % 3329;
                                                                                                                                                                  mul_add_t[0][225] <= (mult_out_1[225] + mult_out_2[225] + mult_out_3[225]) % 3329;
                                                                                                                                                                  mul_add_t[0][226] <= (mult_out_1[226] + mult_out_2[226] + mult_out_3[226]) % 3329;
                                                                                                                                                                  mul_add_t[0][227] <= (mult_out_1[227] + mult_out_2[227] + mult_out_3[227]) % 3329;
                                                                                                                                                                  mul_add_t[0][228] <= (mult_out_1[228] + mult_out_2[228] + mult_out_3[228]) % 3329;
                                                                                                                                                                  mul_add_t[0][229] <= (mult_out_1[229] + mult_out_2[229] + mult_out_3[229]) % 3329;
                                                                                                                                                                  mul_add_t[0][230] <= (mult_out_1[230] + mult_out_2[230] + mult_out_3[230]) % 3329;
                                                                                                                                                                  mul_add_t[0][231] <= (mult_out_1[231] + mult_out_2[231] + mult_out_3[231]) % 3329;
                                                                                                                                                                  mul_add_t[0][232] <= (mult_out_1[232] + mult_out_2[232] + mult_out_3[232]) % 3329;
                                                                                                                                                                  mul_add_t[0][233] <= (mult_out_1[233] + mult_out_2[233] + mult_out_3[233]) % 3329;
                                                                                                                                                                  mul_add_t[0][234] <= (mult_out_1[234] + mult_out_2[234] + mult_out_3[234]) % 3329;
                                                                                                                                                                  mul_add_t[0][235] <= (mult_out_1[235] + mult_out_2[235] + mult_out_3[235]) % 3329;
                                                                                                                                                                  mul_add_t[0][236] <= (mult_out_1[236] + mult_out_2[236] + mult_out_3[236]) % 3329;
                                                                                                                                                                  mul_add_t[0][237] <= (mult_out_1[237] + mult_out_2[237] + mult_out_3[237]) % 3329;
                                                                                                                                                                  mul_add_t[0][238] <= (mult_out_1[238] + mult_out_2[238] + mult_out_3[238]) % 3329;
                                                                                                                                                                  mul_add_t[0][239] <= (mult_out_1[239] + mult_out_2[239] + mult_out_3[239]) % 3329;
                                                                                                                                                                  mul_add_t[0][240] <= (mult_out_1[240] + mult_out_2[240] + mult_out_3[240]) % 3329;
                                                                                                                                                                  mul_add_t[0][241] <= (mult_out_1[241] + mult_out_2[241] + mult_out_3[241]) % 3329;
                                                                                                                                                                  mul_add_t[0][242] <= (mult_out_1[242] + mult_out_2[242] + mult_out_3[242]) % 3329;
                                                                                                                                                                  mul_add_t[0][243] <= (mult_out_1[243] + mult_out_2[243] + mult_out_3[243]) % 3329;
                                                                                                                                                                  mul_add_t[0][244] <= (mult_out_1[244] + mult_out_2[244] + mult_out_3[244]) % 3329;
                                                                                                                                                                  mul_add_t[0][245] <= (mult_out_1[245] + mult_out_2[245] + mult_out_3[245]) % 3329;
                                                                                                                                                                  mul_add_t[0][246] <= (mult_out_1[246] + mult_out_2[246] + mult_out_3[246]) % 3329;
                                                                                                                                                                  mul_add_t[0][247] <= (mult_out_1[247] + mult_out_2[247] + mult_out_3[247]) % 3329;
                                                                                                                                                                  mul_add_t[0][248] <= (mult_out_1[248] + mult_out_2[248] + mult_out_3[248]) % 3329;
                                                                                                                                                                  mul_add_t[0][249] <= (mult_out_1[249] + mult_out_2[249] + mult_out_3[249]) % 3329;
                                                                                                                                                                  mul_add_t[0][250] <= (mult_out_1[250] + mult_out_2[250] + mult_out_3[250]) % 3329;
                                                                                                                                                                  mul_add_t[0][251] <= (mult_out_1[251] + mult_out_2[251] + mult_out_3[251]) % 3329;
                                                                                                                                                                  mul_add_t[0][252] <= (mult_out_1[252] + mult_out_2[252] + mult_out_3[252]) % 3329;
                                                                                                                                                                  mul_add_t[0][253] <= (mult_out_1[253] + mult_out_2[253] + mult_out_3[253]) % 3329;
                                                                                                                                                                  mul_add_t[0][254] <= (mult_out_1[254] + mult_out_2[254] + mult_out_3[254]) % 3329;
                                                                                                                                                                  mul_add_t[0][255] <= (mult_out_1[255] + mult_out_2[255] + mult_out_3[255]) % 3329;
                                                                                                                                                                   mul_add_t[1][0] <= (mult_out_1[0] + mult_out_2[0] + mult_out_3[0]) % 3329;
                                                                                                                                                                         mul_add_t[1][1] <= (mult_out_1[1] + mult_out_2[1] + mult_out_3[1]) % 3329;
                                                                                                                                                                         mul_add_t[1][2] <= (mult_out_1[2] + mult_out_2[2] + mult_out_3[2]) % 3329;
                                                                                                                                                                         mul_add_t[1][3] <= (mult_out_1[3] + mult_out_2[3] + mult_out_3[3]) % 3329;
                                                                                                                                                                         mul_add_t[1][4] <= (mult_out_1[4] + mult_out_2[4] + mult_out_3[4]) % 3329;
                                                                                                                                                                         mul_add_t[1][5] <= (mult_out_1[5] + mult_out_2[5] + mult_out_3[5]) % 3329;
                                                                                                                                                                         mul_add_t[1][6] <= (mult_out_1[6] + mult_out_2[6] + mult_out_3[6]) % 3329;
                                                                                                                                                                         mul_add_t[1][7] <= (mult_out_1[7] + mult_out_2[7] + mult_out_3[7]) % 3329;
                                                                                                                                                                         mul_add_t[1][8] <= (mult_out_1[8] + mult_out_2[8] + mult_out_3[8]) % 3329;
                                                                                                                                                                         mul_add_t[1][9] <= (mult_out_1[9] + mult_out_2[9] + mult_out_3[9]) % 3329;
                                                                                                                                                                         mul_add_t[1][10] <= (mult_out_1[10] + mult_out_2[10] + mult_out_3[10]) % 3329;
                                                                                                                                                                         mul_add_t[1][11] <= (mult_out_1[11] + mult_out_2[11] + mult_out_3[11]) % 3329;
                                                                                                                                                                         mul_add_t[1][12] <= (mult_out_1[12] + mult_out_2[12] + mult_out_3[12]) % 3329;
                                                                                                                                                                         mul_add_t[1][13] <= (mult_out_1[13] + mult_out_2[13] + mult_out_3[13]) % 3329;
                                                                                                                                                                         mul_add_t[1][14] <= (mult_out_1[14] + mult_out_2[14] + mult_out_3[14]) % 3329;
                                                                                                                                                                         mul_add_t[1][15] <= (mult_out_1[15] + mult_out_2[15] + mult_out_3[15]) % 3329;
                                                                                                                                                                         mul_add_t[1][16] <= (mult_out_1[16] + mult_out_2[16] + mult_out_3[16]) % 3329;
                                                                                                                                                                         mul_add_t[1][17] <= (mult_out_1[17] + mult_out_2[17] + mult_out_3[17]) % 3329;
                                                                                                                                                                         mul_add_t[1][18] <= (mult_out_1[18] + mult_out_2[18] + mult_out_3[18]) % 3329;
                                                                                                                                                                         mul_add_t[1][19] <= (mult_out_1[19] + mult_out_2[19] + mult_out_3[19]) % 3329;
                                                                                                                                                                         mul_add_t[1][20] <= (mult_out_1[20] + mult_out_2[20] + mult_out_3[20]) % 3329;
                                                                                                                                                                         mul_add_t[1][21] <= (mult_out_1[21] + mult_out_2[21] + mult_out_3[21]) % 3329;
                                                                                                                                                                         mul_add_t[1][22] <= (mult_out_1[22] + mult_out_2[22] + mult_out_3[22]) % 3329;
                                                                                                                                                                         mul_add_t[1][23] <= (mult_out_1[23] + mult_out_2[23] + mult_out_3[23]) % 3329;
                                                                                                                                                                         mul_add_t[1][24] <= (mult_out_1[24] + mult_out_2[24] + mult_out_3[24]) % 3329;
                                                                                                                                                                         mul_add_t[1][25] <= (mult_out_1[25] + mult_out_2[25] + mult_out_3[25]) % 3329;
                                                                                                                                                                         mul_add_t[1][26] <= (mult_out_1[26] + mult_out_2[26] + mult_out_3[26]) % 3329;
                                                                                                                                                                         mul_add_t[1][27] <= (mult_out_1[27] + mult_out_2[27] + mult_out_3[27]) % 3329;
                                                                                                                                                                         mul_add_t[1][28] <= (mult_out_1[28] + mult_out_2[28] + mult_out_3[28]) % 3329;
                                                                                                                                                                         mul_add_t[1][29] <= (mult_out_1[29] + mult_out_2[29] + mult_out_3[29]) % 3329;
                                                                                                                                                                         mul_add_t[1][30] <= (mult_out_1[30] + mult_out_2[30] + mult_out_3[30]) % 3329;
                                                                                                                                                                         mul_add_t[1][31] <= (mult_out_1[31] + mult_out_2[31] + mult_out_3[31]) % 3329;
                                                                                                                                                                         mul_add_t[1][32] <= (mult_out_1[32] + mult_out_2[32] + mult_out_3[32]) % 3329;
                                                                                                                                                                         mul_add_t[1][33] <= (mult_out_1[33] + mult_out_2[33] + mult_out_3[33]) % 3329;
                                                                                                                                                                         mul_add_t[1][34] <= (mult_out_1[34] + mult_out_2[34] + mult_out_3[34]) % 3329;
                                                                                                                                                                         mul_add_t[1][35] <= (mult_out_1[35] + mult_out_2[35] + mult_out_3[35]) % 3329;
                                                                                                                                                                         mul_add_t[1][36] <= (mult_out_1[36] + mult_out_2[36] + mult_out_3[36]) % 3329;
                                                                                                                                                                         mul_add_t[1][37] <= (mult_out_1[37] + mult_out_2[37] + mult_out_3[37]) % 3329;
                                                                                                                                                                         mul_add_t[1][38] <= (mult_out_1[38] + mult_out_2[38] + mult_out_3[38]) % 3329;
                                                                                                                                                                         mul_add_t[1][39] <= (mult_out_1[39] + mult_out_2[39] + mult_out_3[39]) % 3329;
                                                                                                                                                                         mul_add_t[1][40] <= (mult_out_1[40] + mult_out_2[40] + mult_out_3[40]) % 3329;
                                                                                                                                                                         mul_add_t[1][41] <= (mult_out_1[41] + mult_out_2[41] + mult_out_3[41]) % 3329;
                                                                                                                                                                         mul_add_t[1][42] <= (mult_out_1[42] + mult_out_2[42] + mult_out_3[42]) % 3329;
                                                                                                                                                                         mul_add_t[1][43] <= (mult_out_1[43] + mult_out_2[43] + mult_out_3[43]) % 3329;
                                                                                                                                                                         mul_add_t[1][44] <= (mult_out_1[44] + mult_out_2[44] + mult_out_3[44]) % 3329;
                                                                                                                                                                         mul_add_t[1][45] <= (mult_out_1[45] + mult_out_2[45] + mult_out_3[45]) % 3329;
                                                                                                                                                                         mul_add_t[1][46] <= (mult_out_1[46] + mult_out_2[46] + mult_out_3[46]) % 3329;
                                                                                                                                                                         mul_add_t[1][47] <= (mult_out_1[47] + mult_out_2[47] + mult_out_3[47]) % 3329;
                                                                                                                                                                         mul_add_t[1][48] <= (mult_out_1[48] + mult_out_2[48] + mult_out_3[48]) % 3329;
                                                                                                                                                                         mul_add_t[1][49] <= (mult_out_1[49] + mult_out_2[49] + mult_out_3[49]) % 3329;
                                                                                                                                                                         mul_add_t[1][50] <= (mult_out_1[50] + mult_out_2[50] + mult_out_3[50]) % 3329;
                                                                                                                                                                         mul_add_t[1][51] <= (mult_out_1[51] + mult_out_2[51] + mult_out_3[51]) % 3329;
                                                                                                                                                                         mul_add_t[1][52] <= (mult_out_1[52] + mult_out_2[52] + mult_out_3[52]) % 3329;
                                                                                                                                                                         mul_add_t[1][53] <= (mult_out_1[53] + mult_out_2[53] + mult_out_3[53]) % 3329;
                                                                                                                                                                         mul_add_t[1][54] <= (mult_out_1[54] + mult_out_2[54] + mult_out_3[54]) % 3329;
                                                                                                                                                                         mul_add_t[1][55] <= (mult_out_1[55] + mult_out_2[55] + mult_out_3[55]) % 3329;
                                                                                                                                                                         mul_add_t[1][56] <= (mult_out_1[56] + mult_out_2[56] + mult_out_3[56]) % 3329;
                                                                                                                                                                         mul_add_t[1][57] <= (mult_out_1[57] + mult_out_2[57] + mult_out_3[57]) % 3329;
                                                                                                                                                                         mul_add_t[1][58] <= (mult_out_1[58] + mult_out_2[58] + mult_out_3[58]) % 3329;
                                                                                                                                                                         mul_add_t[1][59] <= (mult_out_1[59] + mult_out_2[59] + mult_out_3[59]) % 3329;
                                                                                                                                                                         mul_add_t[1][60] <= (mult_out_1[60] + mult_out_2[60] + mult_out_3[60]) % 3329;
                                                                                                                                                                         mul_add_t[1][61] <= (mult_out_1[61] + mult_out_2[61] + mult_out_3[61]) % 3329;
                                                                                                                                                                         mul_add_t[1][62] <= (mult_out_1[62] + mult_out_2[62] + mult_out_3[62]) % 3329;
                                                                                                                                                                         mul_add_t[1][63] <= (mult_out_1[63] + mult_out_2[63] + mult_out_3[63]) % 3329;
                                                                                                                                                                         mul_add_t[1][64] <= (mult_out_1[64] + mult_out_2[64] + mult_out_3[64]) % 3329;
                                                                                                                                                                         mul_add_t[1][65] <= (mult_out_1[65] + mult_out_2[65] + mult_out_3[65]) % 3329;
                                                                                                                                                                         mul_add_t[1][66] <= (mult_out_1[66] + mult_out_2[66] + mult_out_3[66]) % 3329;
                                                                                                                                                                         mul_add_t[1][67] <= (mult_out_1[67] + mult_out_2[67] + mult_out_3[67]) % 3329;
                                                                                                                                                                         mul_add_t[1][68] <= (mult_out_1[68] + mult_out_2[68] + mult_out_3[68]) % 3329;
                                                                                                                                                                         mul_add_t[1][69] <= (mult_out_1[69] + mult_out_2[69] + mult_out_3[69]) % 3329;
                                                                                                                                                                         mul_add_t[1][70] <= (mult_out_1[70] + mult_out_2[70] + mult_out_3[70]) % 3329;
                                                                                                                                                                         mul_add_t[1][71] <= (mult_out_1[71] + mult_out_2[71] + mult_out_3[71]) % 3329;
                                                                                                                                                                         mul_add_t[1][72] <= (mult_out_1[72] + mult_out_2[72] + mult_out_3[72]) % 3329;
                                                                                                                                                                         mul_add_t[1][73] <= (mult_out_1[73] + mult_out_2[73] + mult_out_3[73]) % 3329;
                                                                                                                                                                         mul_add_t[1][74] <= (mult_out_1[74] + mult_out_2[74] + mult_out_3[74]) % 3329;
                                                                                                                                                                         mul_add_t[1][75] <= (mult_out_1[75] + mult_out_2[75] + mult_out_3[75]) % 3329;
                                                                                                                                                                         mul_add_t[1][76] <= (mult_out_1[76] + mult_out_2[76] + mult_out_3[76]) % 3329;
                                                                                                                                                                         mul_add_t[1][77] <= (mult_out_1[77] + mult_out_2[77] + mult_out_3[77]) % 3329;
                                                                                                                                                                         mul_add_t[1][78] <= (mult_out_1[78] + mult_out_2[78] + mult_out_3[78]) % 3329;
                                                                                                                                                                         mul_add_t[1][79] <= (mult_out_1[79] + mult_out_2[79] + mult_out_3[79]) % 3329;
                                                                                                                                                                         mul_add_t[1][80] <= (mult_out_1[80] + mult_out_2[80] + mult_out_3[80]) % 3329;
                                                                                                                                                                         mul_add_t[1][81] <= (mult_out_1[81] + mult_out_2[81] + mult_out_3[81]) % 3329;
                                                                                                                                                                         mul_add_t[1][82] <= (mult_out_1[82] + mult_out_2[82] + mult_out_3[82]) % 3329;
                                                                                                                                                                         mul_add_t[1][83] <= (mult_out_1[83] + mult_out_2[83] + mult_out_3[83]) % 3329;
                                                                                                                                                                         mul_add_t[1][84] <= (mult_out_1[84] + mult_out_2[84] + mult_out_3[84]) % 3329;
                                                                                                                                                                         mul_add_t[1][85] <= (mult_out_1[85] + mult_out_2[85] + mult_out_3[85]) % 3329;
                                                                                                                                                                         mul_add_t[1][86] <= (mult_out_1[86] + mult_out_2[86] + mult_out_3[86]) % 3329;
                                                                                                                                                                         mul_add_t[1][87] <= (mult_out_1[87] + mult_out_2[87] + mult_out_3[87]) % 3329;
                                                                                                                                                                         mul_add_t[1][88] <= (mult_out_1[88] + mult_out_2[88] + mult_out_3[88]) % 3329;
                                                                                                                                                                         mul_add_t[1][89] <= (mult_out_1[89] + mult_out_2[89] + mult_out_3[89]) % 3329;
                                                                                                                                                                         mul_add_t[1][90] <= (mult_out_1[90] + mult_out_2[90] + mult_out_3[90]) % 3329;
                                                                                                                                                                         mul_add_t[1][91] <= (mult_out_1[91] + mult_out_2[91] + mult_out_3[91]) % 3329;
                                                                                                                                                                         mul_add_t[1][92] <= (mult_out_1[92] + mult_out_2[92] + mult_out_3[92]) % 3329;
                                                                                                                                                                         mul_add_t[1][93] <= (mult_out_1[93] + mult_out_2[93] + mult_out_3[93]) % 3329;
                                                                                                                                                                         mul_add_t[1][94] <= (mult_out_1[94] + mult_out_2[94] + mult_out_3[94]) % 3329;
                                                                                                                                                                         mul_add_t[1][95] <= (mult_out_1[95] + mult_out_2[95] + mult_out_3[95]) % 3329;
                                                                                                                                                                         mul_add_t[1][96] <= (mult_out_1[96] + mult_out_2[96] + mult_out_3[96]) % 3329;
                                                                                                                                                                         mul_add_t[1][97] <= (mult_out_1[97] + mult_out_2[97] + mult_out_3[97]) % 3329;
                                                                                                                                                                         mul_add_t[1][98] <= (mult_out_1[98] + mult_out_2[98] + mult_out_3[98]) % 3329;
                                                                                                                                                                         mul_add_t[1][99] <= (mult_out_1[99] + mult_out_2[99] + mult_out_3[99]) % 3329;
                                                                                                                                                                         mul_add_t[1][100] <= (mult_out_1[100] + mult_out_2[100] + mult_out_3[100]) % 3329;
                                                                                                                                                                         mul_add_t[1][101] <= (mult_out_1[101] + mult_out_2[101] + mult_out_3[101]) % 3329;
                                                                                                                                                                         mul_add_t[1][102] <= (mult_out_1[102] + mult_out_2[102] + mult_out_3[102]) % 3329;
                                                                                                                                                                         mul_add_t[1][103] <= (mult_out_1[103] + mult_out_2[103] + mult_out_3[103]) % 3329;
                                                                                                                                                                         mul_add_t[1][104] <= (mult_out_1[104] + mult_out_2[104] + mult_out_3[104]) % 3329;
                                                                                                                                                                         mul_add_t[1][105] <= (mult_out_1[105] + mult_out_2[105] + mult_out_3[105]) % 3329;
                                                                                                                                                                         mul_add_t[1][106] <= (mult_out_1[106] + mult_out_2[106] + mult_out_3[106]) % 3329;
                                                                                                                                                                         mul_add_t[1][107] <= (mult_out_1[107] + mult_out_2[107] + mult_out_3[107]) % 3329;
                                                                                                                                                                         mul_add_t[1][108] <= (mult_out_1[108] + mult_out_2[108] + mult_out_3[108]) % 3329;
                                                                                                                                                                         mul_add_t[1][109] <= (mult_out_1[109] + mult_out_2[109] + mult_out_3[109]) % 3329;
                                                                                                                                                                         mul_add_t[1][110] <= (mult_out_1[110] + mult_out_2[110] + mult_out_3[110]) % 3329;
                                                                                                                                                                         mul_add_t[1][111] <= (mult_out_1[111] + mult_out_2[111] + mult_out_3[111]) % 3329;
                                                                                                                                                                         mul_add_t[1][112] <= (mult_out_1[112] + mult_out_2[112] + mult_out_3[112]) % 3329;
                                                                                                                                                                         mul_add_t[1][113] <= (mult_out_1[113] + mult_out_2[113] + mult_out_3[113]) % 3329;
                                                                                                                                                                         mul_add_t[1][114] <= (mult_out_1[114] + mult_out_2[114] + mult_out_3[114]) % 3329;
                                                                                                                                                                         mul_add_t[1][115] <= (mult_out_1[115] + mult_out_2[115] + mult_out_3[115]) % 3329;
                                                                                                                                                                         mul_add_t[1][116] <= (mult_out_1[116] + mult_out_2[116] + mult_out_3[116]) % 3329;
                                                                                                                                                                         mul_add_t[1][117] <= (mult_out_1[117] + mult_out_2[117] + mult_out_3[117]) % 3329;
                                                                                                                                                                         mul_add_t[1][118] <= (mult_out_1[118] + mult_out_2[118] + mult_out_3[118]) % 3329;
                                                                                                                                                                         mul_add_t[1][119] <= (mult_out_1[119] + mult_out_2[119] + mult_out_3[119]) % 3329;
                                                                                                                                                                         mul_add_t[1][120] <= (mult_out_1[120] + mult_out_2[120] + mult_out_3[120]) % 3329;
                                                                                                                                                                         mul_add_t[1][121] <= (mult_out_1[121] + mult_out_2[121] + mult_out_3[121]) % 3329;
                                                                                                                                                                         mul_add_t[1][122] <= (mult_out_1[122] + mult_out_2[122] + mult_out_3[122]) % 3329;
                                                                                                                                                                         mul_add_t[1][123] <= (mult_out_1[123] + mult_out_2[123] + mult_out_3[123]) % 3329;
                                                                                                                                                                         mul_add_t[1][124] <= (mult_out_1[124] + mult_out_2[124] + mult_out_3[124]) % 3329;
                                                                                                                                                                         mul_add_t[1][125] <= (mult_out_1[125] + mult_out_2[125] + mult_out_3[125]) % 3329;
                                                                                                                                                                         mul_add_t[1][126] <= (mult_out_1[126] + mult_out_2[126] + mult_out_3[126]) % 3329;
                                                                                                                                                                         mul_add_t[1][127] <= (mult_out_1[127] + mult_out_2[127] + mult_out_3[127]) % 3329;
                                                                                                                                                                         mul_add_t[1][128] <= (mult_out_1[128] + mult_out_2[128] + mult_out_3[128]) % 3329;
                                                                                                                                                                         mul_add_t[1][129] <= (mult_out_1[129] + mult_out_2[129] + mult_out_3[129]) % 3329;
                                                                                                                                                                         mul_add_t[1][130] <= (mult_out_1[130] + mult_out_2[130] + mult_out_3[130]) % 3329;
                                                                                                                                                                         mul_add_t[1][131] <= (mult_out_1[131] + mult_out_2[131] + mult_out_3[131]) % 3329;
                                                                                                                                                                         mul_add_t[1][132] <= (mult_out_1[132] + mult_out_2[132] + mult_out_3[132]) % 3329;
                                                                                                                                                                         mul_add_t[1][133] <= (mult_out_1[133] + mult_out_2[133] + mult_out_3[133]) % 3329;
                                                                                                                                                                         mul_add_t[1][134] <= (mult_out_1[134] + mult_out_2[134] + mult_out_3[134]) % 3329;
                                                                                                                                                                         mul_add_t[1][135] <= (mult_out_1[135] + mult_out_2[135] + mult_out_3[135]) % 3329;
                                                                                                                                                                         mul_add_t[1][136] <= (mult_out_1[136] + mult_out_2[136] + mult_out_3[136]) % 3329;
                                                                                                                                                                         mul_add_t[1][137] <= (mult_out_1[137] + mult_out_2[137] + mult_out_3[137]) % 3329;
                                                                                                                                                                         mul_add_t[1][138] <= (mult_out_1[138] + mult_out_2[138] + mult_out_3[138]) % 3329;
                                                                                                                                                                         mul_add_t[1][139] <= (mult_out_1[139] + mult_out_2[139] + mult_out_3[139]) % 3329;
                                                                                                                                                                         mul_add_t[1][140] <= (mult_out_1[140] + mult_out_2[140] + mult_out_3[140]) % 3329;
                                                                                                                                                                         mul_add_t[1][141] <= (mult_out_1[141] + mult_out_2[141] + mult_out_3[141]) % 3329;
                                                                                                                                                                         mul_add_t[1][142] <= (mult_out_1[142] + mult_out_2[142] + mult_out_3[142]) % 3329;
                                                                                                                                                                         mul_add_t[1][143] <= (mult_out_1[143] + mult_out_2[143] + mult_out_3[143]) % 3329;
                                                                                                                                                                         mul_add_t[1][144] <= (mult_out_1[144] + mult_out_2[144] + mult_out_3[144]) % 3329;
                                                                                                                                                                         mul_add_t[1][145] <= (mult_out_1[145] + mult_out_2[145] + mult_out_3[145]) % 3329;
                                                                                                                                                                         mul_add_t[1][146] <= (mult_out_1[146] + mult_out_2[146] + mult_out_3[146]) % 3329;
                                                                                                                                                                         mul_add_t[1][147] <= (mult_out_1[147] + mult_out_2[147] + mult_out_3[147]) % 3329;
                                                                                                                                                                         mul_add_t[1][148] <= (mult_out_1[148] + mult_out_2[148] + mult_out_3[148]) % 3329;
                                                                                                                                                                         mul_add_t[1][149] <= (mult_out_1[149] + mult_out_2[149] + mult_out_3[149]) % 3329;
                                                                                                                                                                         mul_add_t[1][150] <= (mult_out_1[150] + mult_out_2[150] + mult_out_3[150]) % 3329;
                                                                                                                                                                         mul_add_t[1][151] <= (mult_out_1[151] + mult_out_2[151] + mult_out_3[151]) % 3329;
                                                                                                                                                                         mul_add_t[1][152] <= (mult_out_1[152] + mult_out_2[152] + mult_out_3[152]) % 3329;
                                                                                                                                                                         mul_add_t[1][153] <= (mult_out_1[153] + mult_out_2[153] + mult_out_3[153]) % 3329;
                                                                                                                                                                         mul_add_t[1][154] <= (mult_out_1[154] + mult_out_2[154] + mult_out_3[154]) % 3329;
                                                                                                                                                                         mul_add_t[1][155] <= (mult_out_1[155] + mult_out_2[155] + mult_out_3[155]) % 3329;
                                                                                                                                                                         mul_add_t[1][156] <= (mult_out_1[156] + mult_out_2[156] + mult_out_3[156]) % 3329;
                                                                                                                                                                         mul_add_t[1][157] <= (mult_out_1[157] + mult_out_2[157] + mult_out_3[157]) % 3329;
                                                                                                                                                                         mul_add_t[1][158] <= (mult_out_1[158] + mult_out_2[158] + mult_out_3[158]) % 3329;
                                                                                                                                                                         mul_add_t[1][159] <= (mult_out_1[159] + mult_out_2[159] + mult_out_3[159]) % 3329;
                                                                                                                                                                         mul_add_t[1][160] <= (mult_out_1[160] + mult_out_2[160] + mult_out_3[160]) % 3329;
                                                                                                                                                                         mul_add_t[1][161] <= (mult_out_1[161] + mult_out_2[161] + mult_out_3[161]) % 3329;
                                                                                                                                                                         mul_add_t[1][162] <= (mult_out_1[162] + mult_out_2[162] + mult_out_3[162]) % 3329;
                                                                                                                                                                         mul_add_t[1][163] <= (mult_out_1[163] + mult_out_2[163] + mult_out_3[163]) % 3329;
                                                                                                                                                                         mul_add_t[1][164] <= (mult_out_1[164] + mult_out_2[164] + mult_out_3[164]) % 3329;
                                                                                                                                                                         mul_add_t[1][165] <= (mult_out_1[165] + mult_out_2[165] + mult_out_3[165]) % 3329;
                                                                                                                                                                         mul_add_t[1][166] <= (mult_out_1[166] + mult_out_2[166] + mult_out_3[166]) % 3329;
                                                                                                                                                                         mul_add_t[1][167] <= (mult_out_1[167] + mult_out_2[167] + mult_out_3[167]) % 3329;
                                                                                                                                                                         mul_add_t[1][168] <= (mult_out_1[168] + mult_out_2[168] + mult_out_3[168]) % 3329;
                                                                                                                                                                         mul_add_t[1][169] <= (mult_out_1[169] + mult_out_2[169] + mult_out_3[169]) % 3329;
                                                                                                                                                                         mul_add_t[1][170] <= (mult_out_1[170] + mult_out_2[170] + mult_out_3[170]) % 3329;
                                                                                                                                                                         mul_add_t[1][171] <= (mult_out_1[171] + mult_out_2[171] + mult_out_3[171]) % 3329;
                                                                                                                                                                         mul_add_t[1][172] <= (mult_out_1[172] + mult_out_2[172] + mult_out_3[172]) % 3329;
                                                                                                                                                                         mul_add_t[1][173] <= (mult_out_1[173] + mult_out_2[173] + mult_out_3[173]) % 3329;
                                                                                                                                                                         mul_add_t[1][174] <= (mult_out_1[174] + mult_out_2[174] + mult_out_3[174]) % 3329;
                                                                                                                                                                         mul_add_t[1][175] <= (mult_out_1[175] + mult_out_2[175] + mult_out_3[175]) % 3329;
                                                                                                                                                                         mul_add_t[1][176] <= (mult_out_1[176] + mult_out_2[176] + mult_out_3[176]) % 3329;
                                                                                                                                                                         mul_add_t[1][177] <= (mult_out_1[177] + mult_out_2[177] + mult_out_3[177]) % 3329;
                                                                                                                                                                         mul_add_t[1][178] <= (mult_out_1[178] + mult_out_2[178] + mult_out_3[178]) % 3329;
                                                                                                                                                                         mul_add_t[1][179] <= (mult_out_1[179] + mult_out_2[179] + mult_out_3[179]) % 3329;
                                                                                                                                                                         mul_add_t[1][180] <= (mult_out_1[180] + mult_out_2[180] + mult_out_3[180]) % 3329;
                                                                                                                                                                         mul_add_t[1][181] <= (mult_out_1[181] + mult_out_2[181] + mult_out_3[181]) % 3329;
                                                                                                                                                                         mul_add_t[1][182] <= (mult_out_1[182] + mult_out_2[182] + mult_out_3[182]) % 3329;
                                                                                                                                                                         mul_add_t[1][183] <= (mult_out_1[183] + mult_out_2[183] + mult_out_3[183]) % 3329;
                                                                                                                                                                         mul_add_t[1][184] <= (mult_out_1[184] + mult_out_2[184] + mult_out_3[184]) % 3329;
                                                                                                                                                                         mul_add_t[1][185] <= (mult_out_1[185] + mult_out_2[185] + mult_out_3[185]) % 3329;
                                                                                                                                                                         mul_add_t[1][186] <= (mult_out_1[186] + mult_out_2[186] + mult_out_3[186]) % 3329;
                                                                                                                                                                         mul_add_t[1][187] <= (mult_out_1[187] + mult_out_2[187] + mult_out_3[187]) % 3329;
                                                                                                                                                                         mul_add_t[1][188] <= (mult_out_1[188] + mult_out_2[188] + mult_out_3[188]) % 3329;
                                                                                                                                                                         mul_add_t[1][189] <= (mult_out_1[189] + mult_out_2[189] + mult_out_3[189]) % 3329;
                                                                                                                                                                         mul_add_t[1][190] <= (mult_out_1[190] + mult_out_2[190] + mult_out_3[190]) % 3329;
                                                                                                                                                                         mul_add_t[1][191] <= (mult_out_1[191] + mult_out_2[191] + mult_out_3[191]) % 3329;
                                                                                                                                                                         mul_add_t[1][192] <= (mult_out_1[192] + mult_out_2[192] + mult_out_3[192]) % 3329;
                                                                                                                                                                         mul_add_t[1][193] <= (mult_out_1[193] + mult_out_2[193] + mult_out_3[193]) % 3329;
                                                                                                                                                                         mul_add_t[1][194] <= (mult_out_1[194] + mult_out_2[194] + mult_out_3[194]) % 3329;
                                                                                                                                                                         mul_add_t[1][195] <= (mult_out_1[195] + mult_out_2[195] + mult_out_3[195]) % 3329;
                                                                                                                                                                         mul_add_t[1][196] <= (mult_out_1[196] + mult_out_2[196] + mult_out_3[196]) % 3329;
                                                                                                                                                                         mul_add_t[1][197] <= (mult_out_1[197] + mult_out_2[197] + mult_out_3[197]) % 3329;
                                                                                                                                                                         mul_add_t[1][198] <= (mult_out_1[198] + mult_out_2[198] + mult_out_3[198]) % 3329;
                                                                                                                                                                         mul_add_t[1][199] <= (mult_out_1[199] + mult_out_2[199] + mult_out_3[199]) % 3329;
                                                                                                                                                                         mul_add_t[1][200] <= (mult_out_1[200] + mult_out_2[200] + mult_out_3[200]) % 3329;
                                                                                                                                                                         mul_add_t[1][201] <= (mult_out_1[201] + mult_out_2[201] + mult_out_3[201]) % 3329;
                                                                                                                                                                         mul_add_t[1][202] <= (mult_out_1[202] + mult_out_2[202] + mult_out_3[202]) % 3329;
                                                                                                                                                                         mul_add_t[1][203] <= (mult_out_1[203] + mult_out_2[203] + mult_out_3[203]) % 3329;
                                                                                                                                                                         mul_add_t[1][204] <= (mult_out_1[204] + mult_out_2[204] + mult_out_3[204]) % 3329;
                                                                                                                                                                         mul_add_t[1][205] <= (mult_out_1[205] + mult_out_2[205] + mult_out_3[205]) % 3329;
                                                                                                                                                                         mul_add_t[1][206] <= (mult_out_1[206] + mult_out_2[206] + mult_out_3[206]) % 3329;
                                                                                                                                                                         mul_add_t[1][207] <= (mult_out_1[207] + mult_out_2[207] + mult_out_3[207]) % 3329;
                                                                                                                                                                         mul_add_t[1][208] <= (mult_out_1[208] + mult_out_2[208] + mult_out_3[208]) % 3329;
                                                                                                                                                                         mul_add_t[1][209] <= (mult_out_1[209] + mult_out_2[209] + mult_out_3[209]) % 3329;
                                                                                                                                                                         mul_add_t[1][210] <= (mult_out_1[210] + mult_out_2[210] + mult_out_3[210]) % 3329;
                                                                                                                                                                         mul_add_t[1][211] <= (mult_out_1[211] + mult_out_2[211] + mult_out_3[211]) % 3329;
                                                                                                                                                                         mul_add_t[1][212] <= (mult_out_1[212] + mult_out_2[212] + mult_out_3[212]) % 3329;
                                                                                                                                                                         mul_add_t[1][213] <= (mult_out_1[213] + mult_out_2[213] + mult_out_3[213]) % 3329;
                                                                                                                                                                         mul_add_t[1][214] <= (mult_out_1[214] + mult_out_2[214] + mult_out_3[214]) % 3329;
                                                                                                                                                                         mul_add_t[1][215] <= (mult_out_1[215] + mult_out_2[215] + mult_out_3[215]) % 3329;
                                                                                                                                                                         mul_add_t[1][216] <= (mult_out_1[216] + mult_out_2[216] + mult_out_3[216]) % 3329;
                                                                                                                                                                         mul_add_t[1][217] <= (mult_out_1[217] + mult_out_2[217] + mult_out_3[217]) % 3329;
                                                                                                                                                                         mul_add_t[1][218] <= (mult_out_1[218] + mult_out_2[218] + mult_out_3[218]) % 3329;
                                                                                                                                                                         mul_add_t[1][219] <= (mult_out_1[219] + mult_out_2[219] + mult_out_3[219]) % 3329;
                                                                                                                                                                         mul_add_t[1][220] <= (mult_out_1[220] + mult_out_2[220] + mult_out_3[220]) % 3329;
                                                                                                                                                                         mul_add_t[1][221] <= (mult_out_1[221] + mult_out_2[221] + mult_out_3[221]) % 3329;
                                                                                                                                                                         mul_add_t[1][222] <= (mult_out_1[222] + mult_out_2[222] + mult_out_3[222]) % 3329;
                                                                                                                                                                         mul_add_t[1][223] <= (mult_out_1[223] + mult_out_2[223] + mult_out_3[223]) % 3329;
                                                                                                                                                                         mul_add_t[1][224] <= (mult_out_1[224] + mult_out_2[224] + mult_out_3[224]) % 3329;
                                                                                                                                                                         mul_add_t[1][225] <= (mult_out_1[225] + mult_out_2[225] + mult_out_3[225]) % 3329;
                                                                                                                                                                         mul_add_t[1][226] <= (mult_out_1[226] + mult_out_2[226] + mult_out_3[226]) % 3329;
                                                                                                                                                                         mul_add_t[1][227] <= (mult_out_1[227] + mult_out_2[227] + mult_out_3[227]) % 3329;
                                                                                                                                                                         mul_add_t[1][228] <= (mult_out_1[228] + mult_out_2[228] + mult_out_3[228]) % 3329;
                                                                                                                                                                         mul_add_t[1][229] <= (mult_out_1[229] + mult_out_2[229] + mult_out_3[229]) % 3329;
                                                                                                                                                                         mul_add_t[1][230] <= (mult_out_1[230] + mult_out_2[230] + mult_out_3[230]) % 3329;
                                                                                                                                                                         mul_add_t[1][231] <= (mult_out_1[231] + mult_out_2[231] + mult_out_3[231]) % 3329;
                                                                                                                                                                         mul_add_t[1][232] <= (mult_out_1[232] + mult_out_2[232] + mult_out_3[232]) % 3329;
                                                                                                                                                                         mul_add_t[1][233] <= (mult_out_1[233] + mult_out_2[233] + mult_out_3[233]) % 3329;
                                                                                                                                                                         mul_add_t[1][234] <= (mult_out_1[234] + mult_out_2[234] + mult_out_3[234]) % 3329;
                                                                                                                                                                         mul_add_t[1][235] <= (mult_out_1[235] + mult_out_2[235] + mult_out_3[235]) % 3329;
                                                                                                                                                                         mul_add_t[1][236] <= (mult_out_1[236] + mult_out_2[236] + mult_out_3[236]) % 3329;
                                                                                                                                                                         mul_add_t[1][237] <= (mult_out_1[237] + mult_out_2[237] + mult_out_3[237]) % 3329;
                                                                                                                                                                         mul_add_t[1][238] <= (mult_out_1[238] + mult_out_2[238] + mult_out_3[238]) % 3329;
                                                                                                                                                                         mul_add_t[1][239] <= (mult_out_1[239] + mult_out_2[239] + mult_out_3[239]) % 3329;
                                                                                                                                                                         mul_add_t[1][240] <= (mult_out_1[240] + mult_out_2[240] + mult_out_3[240]) % 3329;
                                                                                                                                                                         mul_add_t[1][241] <= (mult_out_1[241] + mult_out_2[241] + mult_out_3[241]) % 3329;
                                                                                                                                                                         mul_add_t[1][242] <= (mult_out_1[242] + mult_out_2[242] + mult_out_3[242]) % 3329;
                                                                                                                                                                         mul_add_t[1][243] <= (mult_out_1[243] + mult_out_2[243] + mult_out_3[243]) % 3329;
                                                                                                                                                                         mul_add_t[1][244] <= (mult_out_1[244] + mult_out_2[244] + mult_out_3[244]) % 3329;
                                                                                                                                                                         mul_add_t[1][245] <= (mult_out_1[245] + mult_out_2[245] + mult_out_3[245]) % 3329;
                                                                                                                                                                         mul_add_t[1][246] <= (mult_out_1[246] + mult_out_2[246] + mult_out_3[246]) % 3329;
                                                                                                                                                                         mul_add_t[1][247] <= (mult_out_1[247] + mult_out_2[247] + mult_out_3[247]) % 3329;
                                                                                                                                                                         mul_add_t[1][248] <= (mult_out_1[248] + mult_out_2[248] + mult_out_3[248]) % 3329;
                                                                                                                                                                         mul_add_t[1][249] <= (mult_out_1[249] + mult_out_2[249] + mult_out_3[249]) % 3329;
                                                                                                                                                                         mul_add_t[1][250] <= (mult_out_1[250] + mult_out_2[250] + mult_out_3[250]) % 3329;
                                                                                                                                                                         mul_add_t[1][251] <= (mult_out_1[251] + mult_out_2[251] + mult_out_3[251]) % 3329;
                                                                                                                                                                         mul_add_t[1][252] <= (mult_out_1[252] + mult_out_2[252] + mult_out_3[252]) % 3329;
                                                                                                                                                                         mul_add_t[1][253] <= (mult_out_1[253] + mult_out_2[253] + mult_out_3[253]) % 3329;
                                                                                                                                                                         mul_add_t[1][254] <= (mult_out_1[254] + mult_out_2[254] + mult_out_3[254]) % 3329;
                                                                                                                                                                         mul_add_t[1][255] <= (mult_out_1[255] + mult_out_2[255] + mult_out_3[255]) % 3329;
                                                                                                                                                                         mul_add_t[2][0] <= (mult_out_1[0] + mult_out_2[0] + mult_out_3[0]) % 3329;
                                                                                                                                                                                 mul_add_t[2][1] <= (mult_out_1[1] + mult_out_2[1] + mult_out_3[1]) % 3329;
                                                                                                                                                                                 mul_add_t[2][2] <= (mult_out_1[2] + mult_out_2[2] + mult_out_3[2]) % 3329;
                                                                                                                                                                                 mul_add_t[2][3] <= (mult_out_1[3] + mult_out_2[3] + mult_out_3[3]) % 3329;
                                                                                                                                                                                 mul_add_t[2][4] <= (mult_out_1[4] + mult_out_2[4] + mult_out_3[4]) % 3329;
                                                                                                                                                                                 mul_add_t[2][5] <= (mult_out_1[5] + mult_out_2[5] + mult_out_3[5]) % 3329;
                                                                                                                                                                                 mul_add_t[2][6] <= (mult_out_1[6] + mult_out_2[6] + mult_out_3[6]) % 3329;
                                                                                                                                                                                 mul_add_t[2][7] <= (mult_out_1[7] + mult_out_2[7] + mult_out_3[7]) % 3329;
                                                                                                                                                                                 mul_add_t[2][8] <= (mult_out_1[8] + mult_out_2[8] + mult_out_3[8]) % 3329;
                                                                                                                                                                                 mul_add_t[2][9] <= (mult_out_1[9] + mult_out_2[9] + mult_out_3[9]) % 3329;
                                                                                                                                                                                 mul_add_t[2][10] <= (mult_out_1[10] + mult_out_2[10] + mult_out_3[10]) % 3329;
                                                                                                                                                                                 mul_add_t[2][11] <= (mult_out_1[11] + mult_out_2[11] + mult_out_3[11]) % 3329;
                                                                                                                                                                                 mul_add_t[2][12] <= (mult_out_1[12] + mult_out_2[12] + mult_out_3[12]) % 3329;
                                                                                                                                                                                 mul_add_t[2][13] <= (mult_out_1[13] + mult_out_2[13] + mult_out_3[13]) % 3329;
                                                                                                                                                                                 mul_add_t[2][14] <= (mult_out_1[14] + mult_out_2[14] + mult_out_3[14]) % 3329;
                                                                                                                                                                                 mul_add_t[2][15] <= (mult_out_1[15] + mult_out_2[15] + mult_out_3[15]) % 3329;
                                                                                                                                                                                 mul_add_t[2][16] <= (mult_out_1[16] + mult_out_2[16] + mult_out_3[16]) % 3329;
                                                                                                                                                                                 mul_add_t[2][17] <= (mult_out_1[17] + mult_out_2[17] + mult_out_3[17]) % 3329;
                                                                                                                                                                                 mul_add_t[2][18] <= (mult_out_1[18] + mult_out_2[18] + mult_out_3[18]) % 3329;
                                                                                                                                                                                 mul_add_t[2][19] <= (mult_out_1[19] + mult_out_2[19] + mult_out_3[19]) % 3329;
                                                                                                                                                                                 mul_add_t[2][20] <= (mult_out_1[20] + mult_out_2[20] + mult_out_3[20]) % 3329;
                                                                                                                                                                                 mul_add_t[2][21] <= (mult_out_1[21] + mult_out_2[21] + mult_out_3[21]) % 3329;
                                                                                                                                                                                 mul_add_t[2][22] <= (mult_out_1[22] + mult_out_2[22] + mult_out_3[22]) % 3329;
                                                                                                                                                                                 mul_add_t[2][23] <= (mult_out_1[23] + mult_out_2[23] + mult_out_3[23]) % 3329;
                                                                                                                                                                                 mul_add_t[2][24] <= (mult_out_1[24] + mult_out_2[24] + mult_out_3[24]) % 3329;
                                                                                                                                                                                 mul_add_t[2][25] <= (mult_out_1[25] + mult_out_2[25] + mult_out_3[25]) % 3329;
                                                                                                                                                                                 mul_add_t[2][26] <= (mult_out_1[26] + mult_out_2[26] + mult_out_3[26]) % 3329;
                                                                                                                                                                                 mul_add_t[2][27] <= (mult_out_1[27] + mult_out_2[27] + mult_out_3[27]) % 3329;
                                                                                                                                                                                 mul_add_t[2][28] <= (mult_out_1[28] + mult_out_2[28] + mult_out_3[28]) % 3329;
                                                                                                                                                                                 mul_add_t[2][29] <= (mult_out_1[29] + mult_out_2[29] + mult_out_3[29]) % 3329;
                                                                                                                                                                                 mul_add_t[2][30] <= (mult_out_1[30] + mult_out_2[30] + mult_out_3[30]) % 3329;
                                                                                                                                                                                 mul_add_t[2][31] <= (mult_out_1[31] + mult_out_2[31] + mult_out_3[31]) % 3329;
                                                                                                                                                                                 mul_add_t[2][32] <= (mult_out_1[32] + mult_out_2[32] + mult_out_3[32]) % 3329;
                                                                                                                                                                                 mul_add_t[2][33] <= (mult_out_1[33] + mult_out_2[33] + mult_out_3[33]) % 3329;
                                                                                                                                                                                 mul_add_t[2][34] <= (mult_out_1[34] + mult_out_2[34] + mult_out_3[34]) % 3329;
                                                                                                                                                                                 mul_add_t[2][35] <= (mult_out_1[35] + mult_out_2[35] + mult_out_3[35]) % 3329;
                                                                                                                                                                                 mul_add_t[2][36] <= (mult_out_1[36] + mult_out_2[36] + mult_out_3[36]) % 3329;
                                                                                                                                                                                 mul_add_t[2][37] <= (mult_out_1[37] + mult_out_2[37] + mult_out_3[37]) % 3329;
                                                                                                                                                                                 mul_add_t[2][38] <= (mult_out_1[38] + mult_out_2[38] + mult_out_3[38]) % 3329;
                                                                                                                                                                                 mul_add_t[2][39] <= (mult_out_1[39] + mult_out_2[39] + mult_out_3[39]) % 3329;
                                                                                                                                                                                 mul_add_t[2][40] <= (mult_out_1[40] + mult_out_2[40] + mult_out_3[40]) % 3329;
                                                                                                                                                                                 mul_add_t[2][41] <= (mult_out_1[41] + mult_out_2[41] + mult_out_3[41]) % 3329;
                                                                                                                                                                                 mul_add_t[2][42] <= (mult_out_1[42] + mult_out_2[42] + mult_out_3[42]) % 3329;
                                                                                                                                                                                 mul_add_t[2][43] <= (mult_out_1[43] + mult_out_2[43] + mult_out_3[43]) % 3329;
                                                                                                                                                                                 mul_add_t[2][44] <= (mult_out_1[44] + mult_out_2[44] + mult_out_3[44]) % 3329;
                                                                                                                                                                                 mul_add_t[2][45] <= (mult_out_1[45] + mult_out_2[45] + mult_out_3[45]) % 3329;
                                                                                                                                                                                 mul_add_t[2][46] <= (mult_out_1[46] + mult_out_2[46] + mult_out_3[46]) % 3329;
                                                                                                                                                                                 mul_add_t[2][47] <= (mult_out_1[47] + mult_out_2[47] + mult_out_3[47]) % 3329;
                                                                                                                                                                                 mul_add_t[2][48] <= (mult_out_1[48] + mult_out_2[48] + mult_out_3[48]) % 3329;
                                                                                                                                                                                 mul_add_t[2][49] <= (mult_out_1[49] + mult_out_2[49] + mult_out_3[49]) % 3329;
                                                                                                                                                                                 mul_add_t[2][50] <= (mult_out_1[50] + mult_out_2[50] + mult_out_3[50]) % 3329;
                                                                                                                                                                                 mul_add_t[2][51] <= (mult_out_1[51] + mult_out_2[51] + mult_out_3[51]) % 3329;
                                                                                                                                                                                 mul_add_t[2][52] <= (mult_out_1[52] + mult_out_2[52] + mult_out_3[52]) % 3329;
                                                                                                                                                                                 mul_add_t[2][53] <= (mult_out_1[53] + mult_out_2[53] + mult_out_3[53]) % 3329;
                                                                                                                                                                                 mul_add_t[2][54] <= (mult_out_1[54] + mult_out_2[54] + mult_out_3[54]) % 3329;
                                                                                                                                                                                 mul_add_t[2][55] <= (mult_out_1[55] + mult_out_2[55] + mult_out_3[55]) % 3329;
                                                                                                                                                                                 mul_add_t[2][56] <= (mult_out_1[56] + mult_out_2[56] + mult_out_3[56]) % 3329;
                                                                                                                                                                                 mul_add_t[2][57] <= (mult_out_1[57] + mult_out_2[57] + mult_out_3[57]) % 3329;
                                                                                                                                                                                 mul_add_t[2][58] <= (mult_out_1[58] + mult_out_2[58] + mult_out_3[58]) % 3329;
                                                                                                                                                                                 mul_add_t[2][59] <= (mult_out_1[59] + mult_out_2[59] + mult_out_3[59]) % 3329;
                                                                                                                                                                                 mul_add_t[2][60] <= (mult_out_1[60] + mult_out_2[60] + mult_out_3[60]) % 3329;
                                                                                                                                                                                 mul_add_t[2][61] <= (mult_out_1[61] + mult_out_2[61] + mult_out_3[61]) % 3329;
                                                                                                                                                                                 mul_add_t[2][62] <= (mult_out_1[62] + mult_out_2[62] + mult_out_3[62]) % 3329;
                                                                                                                                                                                 mul_add_t[2][63] <= (mult_out_1[63] + mult_out_2[63] + mult_out_3[63]) % 3329;
                                                                                                                                                                                 mul_add_t[2][64] <= (mult_out_1[64] + mult_out_2[64] + mult_out_3[64]) % 3329;
                                                                                                                                                                                 mul_add_t[2][65] <= (mult_out_1[65] + mult_out_2[65] + mult_out_3[65]) % 3329;
                                                                                                                                                                                 mul_add_t[2][66] <= (mult_out_1[66] + mult_out_2[66] + mult_out_3[66]) % 3329;
                                                                                                                                                                                 mul_add_t[2][67] <= (mult_out_1[67] + mult_out_2[67] + mult_out_3[67]) % 3329;
                                                                                                                                                                                 mul_add_t[2][68] <= (mult_out_1[68] + mult_out_2[68] + mult_out_3[68]) % 3329;
                                                                                                                                                                                 mul_add_t[2][69] <= (mult_out_1[69] + mult_out_2[69] + mult_out_3[69]) % 3329;
                                                                                                                                                                                 mul_add_t[2][70] <= (mult_out_1[70] + mult_out_2[70] + mult_out_3[70]) % 3329;
                                                                                                                                                                                 mul_add_t[2][71] <= (mult_out_1[71] + mult_out_2[71] + mult_out_3[71]) % 3329;
                                                                                                                                                                                 mul_add_t[2][72] <= (mult_out_1[72] + mult_out_2[72] + mult_out_3[72]) % 3329;
                                                                                                                                                                                 mul_add_t[2][73] <= (mult_out_1[73] + mult_out_2[73] + mult_out_3[73]) % 3329;
                                                                                                                                                                                 mul_add_t[2][74] <= (mult_out_1[74] + mult_out_2[74] + mult_out_3[74]) % 3329;
                                                                                                                                                                                 mul_add_t[2][75] <= (mult_out_1[75] + mult_out_2[75] + mult_out_3[75]) % 3329;
                                                                                                                                                                                 mul_add_t[2][76] <= (mult_out_1[76] + mult_out_2[76] + mult_out_3[76]) % 3329;
                                                                                                                                                                                 mul_add_t[2][77] <= (mult_out_1[77] + mult_out_2[77] + mult_out_3[77]) % 3329;
                                                                                                                                                                                 mul_add_t[2][78] <= (mult_out_1[78] + mult_out_2[78] + mult_out_3[78]) % 3329;
                                                                                                                                                                                 mul_add_t[2][79] <= (mult_out_1[79] + mult_out_2[79] + mult_out_3[79]) % 3329;
                                                                                                                                                                                 mul_add_t[2][80] <= (mult_out_1[80] + mult_out_2[80] + mult_out_3[80]) % 3329;
                                                                                                                                                                                 mul_add_t[2][81] <= (mult_out_1[81] + mult_out_2[81] + mult_out_3[81]) % 3329;
                                                                                                                                                                                 mul_add_t[2][82] <= (mult_out_1[82] + mult_out_2[82] + mult_out_3[82]) % 3329;
                                                                                                                                                                                 mul_add_t[2][83] <= (mult_out_1[83] + mult_out_2[83] + mult_out_3[83]) % 3329;
                                                                                                                                                                                 mul_add_t[2][84] <= (mult_out_1[84] + mult_out_2[84] + mult_out_3[84]) % 3329;
                                                                                                                                                                                 mul_add_t[2][85] <= (mult_out_1[85] + mult_out_2[85] + mult_out_3[85]) % 3329;
                                                                                                                                                                                 mul_add_t[2][86] <= (mult_out_1[86] + mult_out_2[86] + mult_out_3[86]) % 3329;
                                                                                                                                                                                 mul_add_t[2][87] <= (mult_out_1[87] + mult_out_2[87] + mult_out_3[87]) % 3329;
                                                                                                                                                                                 mul_add_t[2][88] <= (mult_out_1[88] + mult_out_2[88] + mult_out_3[88]) % 3329;
                                                                                                                                                                                 mul_add_t[2][89] <= (mult_out_1[89] + mult_out_2[89] + mult_out_3[89]) % 3329;
                                                                                                                                                                                 mul_add_t[2][90] <= (mult_out_1[90] + mult_out_2[90] + mult_out_3[90]) % 3329;
                                                                                                                                                                                 mul_add_t[2][91] <= (mult_out_1[91] + mult_out_2[91] + mult_out_3[91]) % 3329;
                                                                                                                                                                                 mul_add_t[2][92] <= (mult_out_1[92] + mult_out_2[92] + mult_out_3[92]) % 3329;
                                                                                                                                                                                 mul_add_t[2][93] <= (mult_out_1[93] + mult_out_2[93] + mult_out_3[93]) % 3329;
                                                                                                                                                                                 mul_add_t[2][94] <= (mult_out_1[94] + mult_out_2[94] + mult_out_3[94]) % 3329;
                                                                                                                                                                                 mul_add_t[2][95] <= (mult_out_1[95] + mult_out_2[95] + mult_out_3[95]) % 3329;
                                                                                                                                                                                 mul_add_t[2][96] <= (mult_out_1[96] + mult_out_2[96] + mult_out_3[96]) % 3329;
                                                                                                                                                                                 mul_add_t[2][97] <= (mult_out_1[97] + mult_out_2[97] + mult_out_3[97]) % 3329;
                                                                                                                                                                                 mul_add_t[2][98] <= (mult_out_1[98] + mult_out_2[98] + mult_out_3[98]) % 3329;
                                                                                                                                                                                 mul_add_t[2][99] <= (mult_out_1[99] + mult_out_2[99] + mult_out_3[99]) % 3329;
                                                                                                                                                                                 mul_add_t[2][100] <= (mult_out_1[100] + mult_out_2[100] + mult_out_3[100]) % 3329;
                                                                                                                                                                                 mul_add_t[2][101] <= (mult_out_1[101] + mult_out_2[101] + mult_out_3[101]) % 3329;
                                                                                                                                                                                 mul_add_t[2][102] <= (mult_out_1[102] + mult_out_2[102] + mult_out_3[102]) % 3329;
                                                                                                                                                                                 mul_add_t[2][103] <= (mult_out_1[103] + mult_out_2[103] + mult_out_3[103]) % 3329;
                                                                                                                                                                                 mul_add_t[2][104] <= (mult_out_1[104] + mult_out_2[104] + mult_out_3[104]) % 3329;
                                                                                                                                                                                 mul_add_t[2][105] <= (mult_out_1[105] + mult_out_2[105] + mult_out_3[105]) % 3329;
                                                                                                                                                                                 mul_add_t[2][106] <= (mult_out_1[106] + mult_out_2[106] + mult_out_3[106]) % 3329;
                                                                                                                                                                                 mul_add_t[2][107] <= (mult_out_1[107] + mult_out_2[107] + mult_out_3[107]) % 3329;
                                                                                                                                                                                 mul_add_t[2][108] <= (mult_out_1[108] + mult_out_2[108] + mult_out_3[108]) % 3329;
                                                                                                                                                                                 mul_add_t[2][109] <= (mult_out_1[109] + mult_out_2[109] + mult_out_3[109]) % 3329;
                                                                                                                                                                                 mul_add_t[2][110] <= (mult_out_1[110] + mult_out_2[110] + mult_out_3[110]) % 3329;
                                                                                                                                                                                 mul_add_t[2][111] <= (mult_out_1[111] + mult_out_2[111] + mult_out_3[111]) % 3329;
                                                                                                                                                                                 mul_add_t[2][112] <= (mult_out_1[112] + mult_out_2[112] + mult_out_3[112]) % 3329;
                                                                                                                                                                                 mul_add_t[2][113] <= (mult_out_1[113] + mult_out_2[113] + mult_out_3[113]) % 3329;
                                                                                                                                                                                 mul_add_t[2][114] <= (mult_out_1[114] + mult_out_2[114] + mult_out_3[114]) % 3329;
                                                                                                                                                                                 mul_add_t[2][115] <= (mult_out_1[115] + mult_out_2[115] + mult_out_3[115]) % 3329;
                                                                                                                                                                                 mul_add_t[2][116] <= (mult_out_1[116] + mult_out_2[116] + mult_out_3[116]) % 3329;
                                                                                                                                                                                 mul_add_t[2][117] <= (mult_out_1[117] + mult_out_2[117] + mult_out_3[117]) % 3329;
                                                                                                                                                                                 mul_add_t[2][118] <= (mult_out_1[118] + mult_out_2[118] + mult_out_3[118]) % 3329;
                                                                                                                                                                                 mul_add_t[2][119] <= (mult_out_1[119] + mult_out_2[119] + mult_out_3[119]) % 3329;
                                                                                                                                                                                 mul_add_t[2][120] <= (mult_out_1[120] + mult_out_2[120] + mult_out_3[120]) % 3329;
                                                                                                                                                                                 mul_add_t[2][121] <= (mult_out_1[121] + mult_out_2[121] + mult_out_3[121]) % 3329;
                                                                                                                                                                                 mul_add_t[2][122] <= (mult_out_1[122] + mult_out_2[122] + mult_out_3[122]) % 3329;
                                                                                                                                                                                 mul_add_t[2][123] <= (mult_out_1[123] + mult_out_2[123] + mult_out_3[123]) % 3329;
                                                                                                                                                                                 mul_add_t[2][124] <= (mult_out_1[124] + mult_out_2[124] + mult_out_3[124]) % 3329;
                                                                                                                                                                                 mul_add_t[2][125] <= (mult_out_1[125] + mult_out_2[125] + mult_out_3[125]) % 3329;
                                                                                                                                                                                 mul_add_t[2][126] <= (mult_out_1[126] + mult_out_2[126] + mult_out_3[126]) % 3329;
                                                                                                                                                                                 mul_add_t[2][127] <= (mult_out_1[127] + mult_out_2[127] + mult_out_3[127]) % 3329;
                                                                                                                                                                                 mul_add_t[2][128] <= (mult_out_1[128] + mult_out_2[128] + mult_out_3[128]) % 3329;
                                                                                                                                                                                 mul_add_t[2][129] <= (mult_out_1[129] + mult_out_2[129] + mult_out_3[129]) % 3329;
                                                                                                                                                                                 mul_add_t[2][130] <= (mult_out_1[130] + mult_out_2[130] + mult_out_3[130]) % 3329;
                                                                                                                                                                                 mul_add_t[2][131] <= (mult_out_1[131] + mult_out_2[131] + mult_out_3[131]) % 3329;
                                                                                                                                                                                 mul_add_t[2][132] <= (mult_out_1[132] + mult_out_2[132] + mult_out_3[132]) % 3329;
                                                                                                                                                                                 mul_add_t[2][133] <= (mult_out_1[133] + mult_out_2[133] + mult_out_3[133]) % 3329;
                                                                                                                                                                                 mul_add_t[2][134] <= (mult_out_1[134] + mult_out_2[134] + mult_out_3[134]) % 3329;
                                                                                                                                                                                 mul_add_t[2][135] <= (mult_out_1[135] + mult_out_2[135] + mult_out_3[135]) % 3329;
                                                                                                                                                                                 mul_add_t[2][136] <= (mult_out_1[136] + mult_out_2[136] + mult_out_3[136]) % 3329;
                                                                                                                                                                                 mul_add_t[2][137] <= (mult_out_1[137] + mult_out_2[137] + mult_out_3[137]) % 3329;
                                                                                                                                                                                 mul_add_t[2][138] <= (mult_out_1[138] + mult_out_2[138] + mult_out_3[138]) % 3329;
                                                                                                                                                                                 mul_add_t[2][139] <= (mult_out_1[139] + mult_out_2[139] + mult_out_3[139]) % 3329;
                                                                                                                                                                                 mul_add_t[2][140] <= (mult_out_1[140] + mult_out_2[140] + mult_out_3[140]) % 3329;
                                                                                                                                                                                 mul_add_t[2][141] <= (mult_out_1[141] + mult_out_2[141] + mult_out_3[141]) % 3329;
                                                                                                                                                                                 mul_add_t[2][142] <= (mult_out_1[142] + mult_out_2[142] + mult_out_3[142]) % 3329;
                                                                                                                                                                                 mul_add_t[2][143] <= (mult_out_1[143] + mult_out_2[143] + mult_out_3[143]) % 3329;
                                                                                                                                                                                 mul_add_t[2][144] <= (mult_out_1[144] + mult_out_2[144] + mult_out_3[144]) % 3329;
                                                                                                                                                                                 mul_add_t[2][145] <= (mult_out_1[145] + mult_out_2[145] + mult_out_3[145]) % 3329;
                                                                                                                                                                                 mul_add_t[2][146] <= (mult_out_1[146] + mult_out_2[146] + mult_out_3[146]) % 3329;
                                                                                                                                                                                 mul_add_t[2][147] <= (mult_out_1[147] + mult_out_2[147] + mult_out_3[147]) % 3329;
                                                                                                                                                                                 mul_add_t[2][148] <= (mult_out_1[148] + mult_out_2[148] + mult_out_3[148]) % 3329;
                                                                                                                                                                                 mul_add_t[2][149] <= (mult_out_1[149] + mult_out_2[149] + mult_out_3[149]) % 3329;
                                                                                                                                                                                 mul_add_t[2][150] <= (mult_out_1[150] + mult_out_2[150] + mult_out_3[150]) % 3329;
                                                                                                                                                                                 mul_add_t[2][151] <= (mult_out_1[151] + mult_out_2[151] + mult_out_3[151]) % 3329;
                                                                                                                                                                                 mul_add_t[2][152] <= (mult_out_1[152] + mult_out_2[152] + mult_out_3[152]) % 3329;
                                                                                                                                                                                 mul_add_t[2][153] <= (mult_out_1[153] + mult_out_2[153] + mult_out_3[153]) % 3329;
                                                                                                                                                                                 mul_add_t[2][154] <= (mult_out_1[154] + mult_out_2[154] + mult_out_3[154]) % 3329;
                                                                                                                                                                                 mul_add_t[2][155] <= (mult_out_1[155] + mult_out_2[155] + mult_out_3[155]) % 3329;
                                                                                                                                                                                 mul_add_t[2][156] <= (mult_out_1[156] + mult_out_2[156] + mult_out_3[156]) % 3329;
                                                                                                                                                                                 mul_add_t[2][157] <= (mult_out_1[157] + mult_out_2[157] + mult_out_3[157]) % 3329;
                                                                                                                                                                                 mul_add_t[2][158] <= (mult_out_1[158] + mult_out_2[158] + mult_out_3[158]) % 3329;
                                                                                                                                                                                 mul_add_t[2][159] <= (mult_out_1[159] + mult_out_2[159] + mult_out_3[159]) % 3329;
                                                                                                                                                                                 mul_add_t[2][160] <= (mult_out_1[160] + mult_out_2[160] + mult_out_3[160]) % 3329;
                                                                                                                                                                                 mul_add_t[2][161] <= (mult_out_1[161] + mult_out_2[161] + mult_out_3[161]) % 3329;
                                                                                                                                                                                 mul_add_t[2][162] <= (mult_out_1[162] + mult_out_2[162] + mult_out_3[162]) % 3329;
                                                                                                                                                                                 mul_add_t[2][163] <= (mult_out_1[163] + mult_out_2[163] + mult_out_3[163]) % 3329;
                                                                                                                                                                                 mul_add_t[2][164] <= (mult_out_1[164] + mult_out_2[164] + mult_out_3[164]) % 3329;
                                                                                                                                                                                 mul_add_t[2][165] <= (mult_out_1[165] + mult_out_2[165] + mult_out_3[165]) % 3329;
                                                                                                                                                                                 mul_add_t[2][166] <= (mult_out_1[166] + mult_out_2[166] + mult_out_3[166]) % 3329;
                                                                                                                                                                                 mul_add_t[2][167] <= (mult_out_1[167] + mult_out_2[167] + mult_out_3[167]) % 3329;
                                                                                                                                                                                 mul_add_t[2][168] <= (mult_out_1[168] + mult_out_2[168] + mult_out_3[168]) % 3329;
                                                                                                                                                                                 mul_add_t[2][169] <= (mult_out_1[169] + mult_out_2[169] + mult_out_3[169]) % 3329;
                                                                                                                                                                                 mul_add_t[2][170] <= (mult_out_1[170] + mult_out_2[170] + mult_out_3[170]) % 3329;
                                                                                                                                                                                 mul_add_t[2][171] <= (mult_out_1[171] + mult_out_2[171] + mult_out_3[171]) % 3329;
                                                                                                                                                                                 mul_add_t[2][172] <= (mult_out_1[172] + mult_out_2[172] + mult_out_3[172]) % 3329;
                                                                                                                                                                                 mul_add_t[2][173] <= (mult_out_1[173] + mult_out_2[173] + mult_out_3[173]) % 3329;
                                                                                                                                                                                 mul_add_t[2][174] <= (mult_out_1[174] + mult_out_2[174] + mult_out_3[174]) % 3329;
                                                                                                                                                                                 mul_add_t[2][175] <= (mult_out_1[175] + mult_out_2[175] + mult_out_3[175]) % 3329;
                                                                                                                                                                                 mul_add_t[2][176] <= (mult_out_1[176] + mult_out_2[176] + mult_out_3[176]) % 3329;
                                                                                                                                                                                 mul_add_t[2][177] <= (mult_out_1[177] + mult_out_2[177] + mult_out_3[177]) % 3329;
                                                                                                                                                                                 mul_add_t[2][178] <= (mult_out_1[178] + mult_out_2[178] + mult_out_3[178]) % 3329;
                                                                                                                                                                                 mul_add_t[2][179] <= (mult_out_1[179] + mult_out_2[179] + mult_out_3[179]) % 3329;
                                                                                                                                                                                 mul_add_t[2][180] <= (mult_out_1[180] + mult_out_2[180] + mult_out_3[180]) % 3329;
                                                                                                                                                                                 mul_add_t[2][181] <= (mult_out_1[181] + mult_out_2[181] + mult_out_3[181]) % 3329;
                                                                                                                                                                                 mul_add_t[2][182] <= (mult_out_1[182] + mult_out_2[182] + mult_out_3[182]) % 3329;
                                                                                                                                                                                 mul_add_t[2][183] <= (mult_out_1[183] + mult_out_2[183] + mult_out_3[183]) % 3329;
                                                                                                                                                                                 mul_add_t[2][184] <= (mult_out_1[184] + mult_out_2[184] + mult_out_3[184]) % 3329;
                                                                                                                                                                                 mul_add_t[2][185] <= (mult_out_1[185] + mult_out_2[185] + mult_out_3[185]) % 3329;
                                                                                                                                                                                 mul_add_t[2][186] <= (mult_out_1[186] + mult_out_2[186] + mult_out_3[186]) % 3329;
                                                                                                                                                                                 mul_add_t[2][187] <= (mult_out_1[187] + mult_out_2[187] + mult_out_3[187]) % 3329;
                                                                                                                                                                                 mul_add_t[2][188] <= (mult_out_1[188] + mult_out_2[188] + mult_out_3[188]) % 3329;
                                                                                                                                                                                 mul_add_t[2][189] <= (mult_out_1[189] + mult_out_2[189] + mult_out_3[189]) % 3329;
                                                                                                                                                                                 mul_add_t[2][190] <= (mult_out_1[190] + mult_out_2[190] + mult_out_3[190]) % 3329;
                                                                                                                                                                                 mul_add_t[2][191] <= (mult_out_1[191] + mult_out_2[191] + mult_out_3[191]) % 3329;
                                                                                                                                                                                 mul_add_t[2][192] <= (mult_out_1[192] + mult_out_2[192] + mult_out_3[192]) % 3329;
                                                                                                                                                                                 mul_add_t[2][193] <= (mult_out_1[193] + mult_out_2[193] + mult_out_3[193]) % 3329;
                                                                                                                                                                                 mul_add_t[2][194] <= (mult_out_1[194] + mult_out_2[194] + mult_out_3[194]) % 3329;
                                                                                                                                                                                 mul_add_t[2][195] <= (mult_out_1[195] + mult_out_2[195] + mult_out_3[195]) % 3329;
                                                                                                                                                                                 mul_add_t[2][196] <= (mult_out_1[196] + mult_out_2[196] + mult_out_3[196]) % 3329;
                                                                                                                                                                                 mul_add_t[2][197] <= (mult_out_1[197] + mult_out_2[197] + mult_out_3[197]) % 3329;
                                                                                                                                                                                 mul_add_t[2][198] <= (mult_out_1[198] + mult_out_2[198] + mult_out_3[198]) % 3329;
                                                                                                                                                                                 mul_add_t[2][199] <= (mult_out_1[199] + mult_out_2[199] + mult_out_3[199]) % 3329;
                                                                                                                                                                                 mul_add_t[2][200] <= (mult_out_1[200] + mult_out_2[200] + mult_out_3[200]) % 3329;
                                                                                                                                                                                 mul_add_t[2][201] <= (mult_out_1[201] + mult_out_2[201] + mult_out_3[201]) % 3329;
                                                                                                                                                                                 mul_add_t[2][202] <= (mult_out_1[202] + mult_out_2[202] + mult_out_3[202]) % 3329;
                                                                                                                                                                                 mul_add_t[2][203] <= (mult_out_1[203] + mult_out_2[203] + mult_out_3[203]) % 3329;
                                                                                                                                                                                 mul_add_t[2][204] <= (mult_out_1[204] + mult_out_2[204] + mult_out_3[204]) % 3329;
                                                                                                                                                                                 mul_add_t[2][205] <= (mult_out_1[205] + mult_out_2[205] + mult_out_3[205]) % 3329;
                                                                                                                                                                                 mul_add_t[2][206] <= (mult_out_1[206] + mult_out_2[206] + mult_out_3[206]) % 3329;
                                                                                                                                                                                 mul_add_t[2][207] <= (mult_out_1[207] + mult_out_2[207] + mult_out_3[207]) % 3329;
                                                                                                                                                                                 mul_add_t[2][208] <= (mult_out_1[208] + mult_out_2[208] + mult_out_3[208]) % 3329;
                                                                                                                                                                                 mul_add_t[2][209] <= (mult_out_1[209] + mult_out_2[209] + mult_out_3[209]) % 3329;
                                                                                                                                                                                 mul_add_t[2][210] <= (mult_out_1[210] + mult_out_2[210] + mult_out_3[210]) % 3329;
                                                                                                                                                                                 mul_add_t[2][211] <= (mult_out_1[211] + mult_out_2[211] + mult_out_3[211]) % 3329;
                                                                                                                                                                                 mul_add_t[2][212] <= (mult_out_1[212] + mult_out_2[212] + mult_out_3[212]) % 3329;
                                                                                                                                                                                 mul_add_t[2][213] <= (mult_out_1[213] + mult_out_2[213] + mult_out_3[213]) % 3329;
                                                                                                                                                                                 mul_add_t[2][214] <= (mult_out_1[214] + mult_out_2[214] + mult_out_3[214]) % 3329;
                                                                                                                                                                                 mul_add_t[2][215] <= (mult_out_1[215] + mult_out_2[215] + mult_out_3[215]) % 3329;
                                                                                                                                                                                 mul_add_t[2][216] <= (mult_out_1[216] + mult_out_2[216] + mult_out_3[216]) % 3329;
                                                                                                                                                                                 mul_add_t[2][217] <= (mult_out_1[217] + mult_out_2[217] + mult_out_3[217]) % 3329;
                                                                                                                                                                                 mul_add_t[2][218] <= (mult_out_1[218] + mult_out_2[218] + mult_out_3[218]) % 3329;
                                                                                                                                                                                 mul_add_t[2][219] <= (mult_out_1[219] + mult_out_2[219] + mult_out_3[219]) % 3329;
                                                                                                                                                                                 mul_add_t[2][220] <= (mult_out_1[220] + mult_out_2[220] + mult_out_3[220]) % 3329;
                                                                                                                                                                                 mul_add_t[2][221] <= (mult_out_1[221] + mult_out_2[221] + mult_out_3[221]) % 3329;
                                                                                                                                                                                 mul_add_t[2][222] <= (mult_out_1[222] + mult_out_2[222] + mult_out_3[222]) % 3329;
                                                                                                                                                                                 mul_add_t[2][223] <= (mult_out_1[223] + mult_out_2[223] + mult_out_3[223]) % 3329;
                                                                                                                                                                                 mul_add_t[2][224] <= (mult_out_1[224] + mult_out_2[224] + mult_out_3[224]) % 3329;
                                                                                                                                                                                 mul_add_t[2][225] <= (mult_out_1[225] + mult_out_2[225] + mult_out_3[225]) % 3329;
                                                                                                                                                                                 mul_add_t[2][226] <= (mult_out_1[226] + mult_out_2[226] + mult_out_3[226]) % 3329;
                                                                                                                                                                                 mul_add_t[2][227] <= (mult_out_1[227] + mult_out_2[227] + mult_out_3[227]) % 3329;
                                                                                                                                                                                 mul_add_t[2][228] <= (mult_out_1[228] + mult_out_2[228] + mult_out_3[228]) % 3329;
                                                                                                                                                                                 mul_add_t[2][229] <= (mult_out_1[229] + mult_out_2[229] + mult_out_3[229]) % 3329;
                                                                                                                                                                                 mul_add_t[2][230] <= (mult_out_1[230] + mult_out_2[230] + mult_out_3[230]) % 3329;
                                                                                                                                                                                 mul_add_t[2][231] <= (mult_out_1[231] + mult_out_2[231] + mult_out_3[231]) % 3329;
                                                                                                                                                                                 mul_add_t[2][232] <= (mult_out_1[232] + mult_out_2[232] + mult_out_3[232]) % 3329;
                                                                                                                                                                                 mul_add_t[2][233] <= (mult_out_1[233] + mult_out_2[233] + mult_out_3[233]) % 3329;
                                                                                                                                                                                 mul_add_t[2][234] <= (mult_out_1[234] + mult_out_2[234] + mult_out_3[234]) % 3329;
                                                                                                                                                                                 mul_add_t[2][235] <= (mult_out_1[235] + mult_out_2[235] + mult_out_3[235]) % 3329;
                                                                                                                                                                                 mul_add_t[2][236] <= (mult_out_1[236] + mult_out_2[236] + mult_out_3[236]) % 3329;
                                                                                                                                                                                 mul_add_t[2][237] <= (mult_out_1[237] + mult_out_2[237] + mult_out_3[237]) % 3329;
                                                                                                                                                                                 mul_add_t[2][238] <= (mult_out_1[238] + mult_out_2[238] + mult_out_3[238]) % 3329;
                                                                                                                                                                                 mul_add_t[2][239] <= (mult_out_1[239] + mult_out_2[239] + mult_out_3[239]) % 3329;
                                                                                                                                                                                 mul_add_t[2][240] <= (mult_out_1[240] + mult_out_2[240] + mult_out_3[240]) % 3329;
                                                                                                                                                                                 mul_add_t[2][241] <= (mult_out_1[241] + mult_out_2[241] + mult_out_3[241]) % 3329;
                                                                                                                                                                                 mul_add_t[2][242] <= (mult_out_1[242] + mult_out_2[242] + mult_out_3[242]) % 3329;
                                                                                                                                                                                 mul_add_t[2][243] <= (mult_out_1[243] + mult_out_2[243] + mult_out_3[243]) % 3329;
                                                                                                                                                                                 mul_add_t[2][244] <= (mult_out_1[244] + mult_out_2[244] + mult_out_3[244]) % 3329;
                                                                                                                                                                                 mul_add_t[2][245] <= (mult_out_1[245] + mult_out_2[245] + mult_out_3[245]) % 3329;
                                                                                                                                                                                 mul_add_t[2][246] <= (mult_out_1[246] + mult_out_2[246] + mult_out_3[246]) % 3329;
                                                                                                                                                                                 mul_add_t[2][247] <= (mult_out_1[247] + mult_out_2[247] + mult_out_3[247]) % 3329;
                                                                                                                                                                                 mul_add_t[2][248] <= (mult_out_1[248] + mult_out_2[248] + mult_out_3[248]) % 3329;
                                                                                                                                                                                 mul_add_t[2][249] <= (mult_out_1[249] + mult_out_2[249] + mult_out_3[249]) % 3329;
                                                                                                                                                                                 mul_add_t[2][250] <= (mult_out_1[250] + mult_out_2[250] + mult_out_3[250]) % 3329;
                                                                                                                                                                                 mul_add_t[2][251] <= (mult_out_1[251] + mult_out_2[251] + mult_out_3[251]) % 3329;
                                                                                                                                                                                 mul_add_t[2][252] <= (mult_out_1[252] + mult_out_2[252] + mult_out_3[252]) % 3329;
                                                                                                                                                                                 mul_add_t[2][253] <= (mult_out_1[253] + mult_out_2[253] + mult_out_3[253]) % 3329;
                                                                                                                                                                                 mul_add_t[2][254] <= (mult_out_1[254] + mult_out_2[254] + mult_out_3[254]) % 3329;
                                                                                                                                                                                 mul_add_t[2][255] <= (mult_out_1[255] + mult_out_2[255] + mult_out_3[255]) % 3329;
                                                                                                                                                                                 u[0][0] = in_1[0] + e1[0][0] %3329;
                                                                                                                                                                                 u[0][1] = in_1[1] + e1[0][1] %3329;
                                                                                                                                                                                 u[0][2] = in_1[2] + e1[0][2] %3329;
                                                                                                                                                                                 u[0][3] = in_1[3] + e1[0][3] %3329;
                                                                                                                                                                                 u[0][4] = in_1[4] + e1[0][4] %3329;
                                                                                                                                                                                 u[0][5] = in_1[5] + e1[0][5] %3329;
                                                                                                                                                                                 u[0][6] = in_1[6] + e1[0][6] %3329;
                                                                                                                                                                                 u[0][7] = in_1[7] + e1[0][7] %3329;
                                                                                                                                                                                 u[0][8] = in_1[8] + e1[0][8] %3329;
                                                                                                                                                                                 u[0][9] = in_1[9] + e1[0][9] %3329;
                                                                                                                                                                                 u[0][10] = in_1[10] + e1[0][10] %3329;
                                                                                                                                                                                 u[0][11] = in_1[11] + e1[0][11] %3329;
                                                                                                                                                                                 u[0][12] = in_1[12] + e1[0][12] %3329;
                                                                                                                                                                                 u[0][13] = in_1[13] + e1[0][13] %3329;
                                                                                                                                                                                 u[0][14] = in_1[14] + e1[0][14] %3329;
                                                                                                                                                                                 u[0][15] = in_1[15] + e1[0][15] %3329;
                                                                                                                                                                                 u[0][16] = in_1[16] + e1[0][16] %3329;
                                                                                                                                                                                 u[0][17] = in_1[17] + e1[0][17] %3329;
                                                                                                                                                                                 u[0][18] = in_1[18] + e1[0][18] %3329;
                                                                                                                                                                                 u[0][19] = in_1[19] + e1[0][19] %3329;
                                                                                                                                                                                 u[0][20] = in_1[20] + e1[0][20] %3329;
                                                                                                                                                                                 u[0][21] = in_1[21] + e1[0][21] %3329;
                                                                                                                                                                                 u[0][22] = in_1[22] + e1[0][22] %3329;
                                                                                                                                                                                 u[0][23] = in_1[23] + e1[0][23] %3329;
                                                                                                                                                                                 u[0][24] = in_1[24] + e1[0][24] %3329;
                                                                                                                                                                                 u[0][25] = in_1[25] + e1[0][25] %3329;
                                                                                                                                                                                 u[0][26] = in_1[26] + e1[0][26] %3329;
                                                                                                                                                                                 u[0][27] = in_1[27] + e1[0][27] %3329;
                                                                                                                                                                                 u[0][28] = in_1[28] + e1[0][28] %3329;
                                                                                                                                                                                 u[0][29] = in_1[29] + e1[0][29] %3329;
                                                                                                                                                                                 u[0][30] = in_1[30] + e1[0][30] %3329;
                                                                                                                                                                                 u[0][31] = in_1[31] + e1[0][31] %3329;
                                                                                                                                                                                 u[0][32] = in_1[32] + e1[0][32] %3329;
                                                                                                                                                                                 u[0][33] = in_1[33] + e1[0][33] %3329;
                                                                                                                                                                                 u[0][34] = in_1[34] + e1[0][34] %3329;
                                                                                                                                                                                 u[0][35] = in_1[35] + e1[0][35] %3329;
                                                                                                                                                                                 u[0][36] = in_1[36] + e1[0][36] %3329;
                                                                                                                                                                                 u[0][37] = in_1[37] + e1[0][37] %3329;
                                                                                                                                                                                 u[0][38] = in_1[38] + e1[0][38] %3329;
                                                                                                                                                                                 u[0][39] = in_1[39] + e1[0][39] %3329;
                                                                                                                                                                                 u[0][40] = in_1[40] + e1[0][40] %3329;
                                                                                                                                                                                 u[0][41] = in_1[41] + e1[0][41] %3329;
                                                                                                                                                                                 u[0][42] = in_1[42] + e1[0][42] %3329;
                                                                                                                                                                                 u[0][43] = in_1[43] + e1[0][43] %3329;
                                                                                                                                                                                 u[0][44] = in_1[44] + e1[0][44] %3329;
                                                                                                                                                                                 u[0][45] = in_1[45] + e1[0][45] %3329;
                                                                                                                                                                                 u[0][46] = in_1[46] + e1[0][46] %3329;
                                                                                                                                                                                 u[0][47] = in_1[47] + e1[0][47] %3329;
                                                                                                                                                                                 u[0][48] = in_1[48] + e1[0][48] %3329;
                                                                                                                                                                                 u[0][49] = in_1[49] + e1[0][49] %3329;
                                                                                                                                                                                 u[0][50] = in_1[50] + e1[0][50] %3329;
                                                                                                                                                                                 u[0][51] = in_1[51] + e1[0][51] %3329;
                                                                                                                                                                                 u[0][52] = in_1[52] + e1[0][52] %3329;
                                                                                                                                                                                 u[0][53] = in_1[53] + e1[0][53] %3329;
                                                                                                                                                                                 u[0][54] = in_1[54] + e1[0][54] %3329;
                                                                                                                                                                                 u[0][55] = in_1[55] + e1[0][55] %3329;
                                                                                                                                                                                 u[0][56] = in_1[56] + e1[0][56] %3329;
                                                                                                                                                                                 u[0][57] = in_1[57] + e1[0][57] %3329;
                                                                                                                                                                                 u[0][58] = in_1[58] + e1[0][58] %3329;
                                                                                                                                                                                 u[0][59] = in_1[59] + e1[0][59] %3329;
                                                                                                                                                                                 u[0][60] = in_1[60] + e1[0][60] %3329;
                                                                                                                                                                                 u[0][61] = in_1[61] + e1[0][61] %3329;
                                                                                                                                                                                 u[0][62] = in_1[62] + e1[0][62] %3329;
                                                                                                                                                                                 u[0][63] = in_1[63] + e1[0][63] %3329;
                                                                                                                                                                                 u[0][64] = in_1[64] + e1[0][64] %3329;
                                                                                                                                                                                 u[0][65] = in_1[65] + e1[0][65] %3329;
                                                                                                                                                                                 u[0][66] = in_1[66] + e1[0][66] %3329;
                                                                                                                                                                                 u[0][67] = in_1[67] + e1[0][67] %3329;
                                                                                                                                                                                 u[0][68] = in_1[68] + e1[0][68] %3329;
                                                                                                                                                                                 u[0][69] = in_1[69] + e1[0][69] %3329;
                                                                                                                                                                                 u[0][70] = in_1[70] + e1[0][70] %3329;
                                                                                                                                                                                 u[0][71] = in_1[71] + e1[0][71] %3329;
                                                                                                                                                                                 u[0][72] = in_1[72] + e1[0][72] %3329;
                                                                                                                                                                                 u[0][73] = in_1[73] + e1[0][73] %3329;
                                                                                                                                                                                 u[0][74] = in_1[74] + e1[0][74] %3329;
                                                                                                                                                                                 u[0][75] = in_1[75] + e1[0][75] %3329;
                                                                                                                                                                                 u[0][76] = in_1[76] + e1[0][76] %3329;
                                                                                                                                                                                 u[0][77] = in_1[77] + e1[0][77] %3329;
                                                                                                                                                                                 u[0][78] = in_1[78] + e1[0][78] %3329;
                                                                                                                                                                                 u[0][79] = in_1[79] + e1[0][79] %3329;
                                                                                                                                                                                 u[0][80] = in_1[80] + e1[0][80] %3329;
                                                                                                                                                                                 u[0][81] = in_1[81] + e1[0][81] %3329;
                                                                                                                                                                                 u[0][82] = in_1[82] + e1[0][82] %3329;
                                                                                                                                                                                 u[0][83] = in_1[83] + e1[0][83] %3329;
                                                                                                                                                                                 u[0][84] = in_1[84] + e1[0][84] %3329;
                                                                                                                                                                                 u[0][85] = in_1[85] + e1[0][85] %3329;
                                                                                                                                                                                 u[0][86] = in_1[86] + e1[0][86] %3329;
                                                                                                                                                                                 u[0][87] = in_1[87] + e1[0][87] %3329;
                                                                                                                                                                                 u[0][88] = in_1[88] + e1[0][88] %3329;
                                                                                                                                                                                 u[0][89] = in_1[89] + e1[0][89] %3329;
                                                                                                                                                                                 u[0][90] = in_1[90] + e1[0][90] %3329;
                                                                                                                                                                                 u[0][91] = in_1[91] + e1[0][91] %3329;
                                                                                                                                                                                 u[0][92] = in_1[92] + e1[0][92] %3329;
                                                                                                                                                                                 u[0][93] = in_1[93] + e1[0][93] %3329;
                                                                                                                                                                                 u[0][94] = in_1[94] + e1[0][94] %3329;
                                                                                                                                                                                 u[0][95] = in_1[95] + e1[0][95] %3329;
                                                                                                                                                                                 u[0][96] = in_1[96] + e1[0][96] %3329;
                                                                                                                                                                                 u[0][97] = in_1[97] + e1[0][97] %3329;
                                                                                                                                                                                 u[0][98] = in_1[98] + e1[0][98] %3329;
                                                                                                                                                                                 u[0][99] = in_1[99] + e1[0][99] %3329;
                                                                                                                                                                                 u[0][100] = in_1[100] + e1[0][100] %3329;
                                                                                                                                                                                 u[0][101] = in_1[101] + e1[0][101] %3329;
                                                                                                                                                                                 u[0][102] = in_1[102] + e1[0][102] %3329;
                                                                                                                                                                                 u[0][103] = in_1[103] + e1[0][103] %3329;
                                                                                                                                                                                 u[0][104] = in_1[104] + e1[0][104] %3329;
                                                                                                                                                                                 u[0][105] = in_1[105] + e1[0][105] %3329;
                                                                                                                                                                                 u[0][106] = in_1[106] + e1[0][106] %3329;
                                                                                                                                                                                 u[0][107] = in_1[107] + e1[0][107] %3329;
                                                                                                                                                                                 u[0][108] = in_1[108] + e1[0][108] %3329;
                                                                                                                                                                                 u[0][109] = in_1[109] + e1[0][109] %3329;
                                                                                                                                                                                 u[0][110] = in_1[110] + e1[0][110] %3329;
                                                                                                                                                                                 u[0][111] = in_1[111] + e1[0][111] %3329;
                                                                                                                                                                                 u[0][112] = in_1[112] + e1[0][112] %3329;
                                                                                                                                                                                 u[0][113] = in_1[113] + e1[0][113] %3329;
                                                                                                                                                                                 u[0][114] = in_1[114] + e1[0][114] %3329;
                                                                                                                                                                                 u[0][115] = in_1[115] + e1[0][115] %3329;
                                                                                                                                                                                 u[0][116] = in_1[116] + e1[0][116] %3329;
                                                                                                                                                                                 u[0][117] = in_1[117] + e1[0][117] %3329;
                                                                                                                                                                                 u[0][118] = in_1[118] + e1[0][118] %3329;
                                                                                                                                                                                 u[0][119] = in_1[119] + e1[0][119] %3329;
                                                                                                                                                                                 u[0][120] = in_1[120] + e1[0][120] %3329;
                                                                                                                                                                                 u[0][121] = in_1[121] + e1[0][121] %3329;
                                                                                                                                                                                 u[0][122] = in_1[122] + e1[0][122] %3329;
                                                                                                                                                                                 u[0][123] = in_1[123] + e1[0][123] %3329;
                                                                                                                                                                                 u[0][124] = in_1[124] + e1[0][124] %3329;
                                                                                                                                                                                 u[0][125] = in_1[125] + e1[0][125] %3329;
                                                                                                                                                                                 u[0][126] = in_1[126] + e1[0][126] %3329;
                                                                                                                                                                                 u[0][127] = in_1[127] + e1[0][127] %3329;
                                                                                                                                                                                 u[0][128] = in_1[128] + e1[0][128] %3329;
                                                                                                                                                                                 u[0][129] = in_1[129] + e1[0][129] %3329;
                                                                                                                                                                                 u[0][130] = in_1[130] + e1[0][130] %3329;
                                                                                                                                                                                 u[0][131] = in_1[131] + e1[0][131] %3329;
                                                                                                                                                                                 u[0][132] = in_1[132] + e1[0][132] %3329;
                                                                                                                                                                                 u[0][133] = in_1[133] + e1[0][133] %3329;
                                                                                                                                                                                 u[0][134] = in_1[134] + e1[0][134] %3329;
                                                                                                                                                                                 u[0][135] = in_1[135] + e1[0][135] %3329;
                                                                                                                                                                                 u[0][136] = in_1[136] + e1[0][136] %3329;
                                                                                                                                                                                 u[0][137] = in_1[137] + e1[0][137] %3329;
                                                                                                                                                                                 u[0][138] = in_1[138] + e1[0][138] %3329;
                                                                                                                                                                                 u[0][139] = in_1[139] + e1[0][139] %3329;
                                                                                                                                                                                 u[0][140] = in_1[140] + e1[0][140] %3329;
                                                                                                                                                                                 u[0][141] = in_1[141] + e1[0][141] %3329;
                                                                                                                                                                                 u[0][142] = in_1[142] + e1[0][142] %3329;
                                                                                                                                                                                 u[0][143] = in_1[143] + e1[0][143] %3329;
                                                                                                                                                                                 u[0][144] = in_1[144] + e1[0][144] %3329;
                                                                                                                                                                                 u[0][145] = in_1[145] + e1[0][145] %3329;
                                                                                                                                                                                 u[0][146] = in_1[146] + e1[0][146] %3329;
                                                                                                                                                                                 u[0][147] = in_1[147] + e1[0][147] %3329;
                                                                                                                                                                                 u[0][148] = in_1[148] + e1[0][148] %3329;
                                                                                                                                                                                 u[0][149] = in_1[149] + e1[0][149] %3329;
                                                                                                                                                                                 u[0][150] = in_1[150] + e1[0][150] %3329;
                                                                                                                                                                                 u[0][151] = in_1[151] + e1[0][151] %3329;
                                                                                                                                                                                 u[0][152] = in_1[152] + e1[0][152] %3329;
                                                                                                                                                                                 u[0][153] = in_1[153] + e1[0][153] %3329;
                                                                                                                                                                                 u[0][154] = in_1[154] + e1[0][154] %3329;
                                                                                                                                                                                 u[0][155] = in_1[155] + e1[0][155] %3329;
                                                                                                                                                                                 u[0][156] = in_1[156] + e1[0][156] %3329;
                                                                                                                                                                                 u[0][157] = in_1[157] + e1[0][157] %3329;
                                                                                                                                                                                 u[0][158] = in_1[158] + e1[0][158] %3329;
                                                                                                                                                                                 u[0][159] = in_1[159] + e1[0][159] %3329;
                                                                                                                                                                                 u[0][160] = in_1[160] + e1[0][160] %3329;
                                                                                                                                                                                 u[0][161] = in_1[161] + e1[0][161] %3329;
                                                                                                                                                                                 u[0][162] = in_1[162] + e1[0][162] %3329;
                                                                                                                                                                                 u[0][163] = in_1[163] + e1[0][163] %3329;
                                                                                                                                                                                 u[0][164] = in_1[164] + e1[0][164] %3329;
                                                                                                                                                                                 u[0][165] = in_1[165] + e1[0][165] %3329;
                                                                                                                                                                                 u[0][166] = in_1[166] + e1[0][166] %3329;
                                                                                                                                                                                 u[0][167] = in_1[167] + e1[0][167] %3329;
                                                                                                                                                                                 u[0][168] = in_1[168] + e1[0][168] %3329;
                                                                                                                                                                                 u[0][169] = in_1[169] + e1[0][169] %3329;
                                                                                                                                                                                 u[0][170] = in_1[170] + e1[0][170] %3329;
                                                                                                                                                                                 u[0][171] = in_1[171] + e1[0][171] %3329;
                                                                                                                                                                                 u[0][172] = in_1[172] + e1[0][172] %3329;
                                                                                                                                                                                 u[0][173] = in_1[173] + e1[0][173] %3329;
                                                                                                                                                                                 u[0][174] = in_1[174] + e1[0][174] %3329;
                                                                                                                                                                                 u[0][175] = in_1[175] + e1[0][175] %3329;
                                                                                                                                                                                 u[0][176] = in_1[176] + e1[0][176] %3329;
                                                                                                                                                                                 u[0][177] = in_1[177] + e1[0][177] %3329;
                                                                                                                                                                                 u[0][178] = in_1[178] + e1[0][178] %3329;
                                                                                                                                                                                 u[0][179] = in_1[179] + e1[0][179] %3329;
                                                                                                                                                                                 u[0][180] = in_1[180] + e1[0][180] %3329;
                                                                                                                                                                                 u[0][181] = in_1[181] + e1[0][181] %3329;
                                                                                                                                                                                 u[0][182] = in_1[182] + e1[0][182] %3329;
                                                                                                                                                                                 u[0][183] = in_1[183] + e1[0][183] %3329;
                                                                                                                                                                                 u[0][184] = in_1[184] + e1[0][184] %3329;
                                                                                                                                                                                 u[0][185] = in_1[185] + e1[0][185] %3329;
                                                                                                                                                                                 u[0][186] = in_1[186] + e1[0][186] %3329;
                                                                                                                                                                                 u[0][187] = in_1[187] + e1[0][187] %3329;
                                                                                                                                                                                 u[0][188] = in_1[188] + e1[0][188] %3329;
                                                                                                                                                                                 u[0][189] = in_1[189] + e1[0][189] %3329;
                                                                                                                                                                                 u[0][190] = in_1[190] + e1[0][190] %3329;
                                                                                                                                                                                 u[0][191] = in_1[191] + e1[0][191] %3329;
                                                                                                                                                                                 u[0][192] = in_1[192] + e1[0][192] %3329;
                                                                                                                                                                                 u[0][193] = in_1[193] + e1[0][193] %3329;
                                                                                                                                                                                 u[0][194] = in_1[194] + e1[0][194] %3329;
                                                                                                                                                                                 u[0][195] = in_1[195] + e1[0][195] %3329;
                                                                                                                                                                                 u[0][196] = in_1[196] + e1[0][196] %3329;
                                                                                                                                                                                 u[0][197] = in_1[197] + e1[0][197] %3329;
                                                                                                                                                                                 u[0][198] = in_1[198] + e1[0][198] %3329;
                                                                                                                                                                                 u[0][199] = in_1[199] + e1[0][199] %3329;
                                                                                                                                                                                 u[0][200] = in_1[200] + e1[0][200] %3329;
                                                                                                                                                                                 u[0][201] = in_1[201] + e1[0][201] %3329;
                                                                                                                                                                                 u[0][202] = in_1[202] + e1[0][202] %3329;
                                                                                                                                                                                 u[0][203] = in_1[203] + e1[0][203] %3329;
                                                                                                                                                                                 u[0][204] = in_1[204] + e1[0][204] %3329;
                                                                                                                                                                                 u[0][205] = in_1[205] + e1[0][205] %3329;
                                                                                                                                                                                 u[0][206] = in_1[206] + e1[0][206] %3329;
                                                                                                                                                                                 u[0][207] = in_1[207] + e1[0][207] %3329;
                                                                                                                                                                                 u[0][208] = in_1[208] + e1[0][208] %3329;
                                                                                                                                                                                 u[0][209] = in_1[209] + e1[0][209] %3329;
                                                                                                                                                                                 u[0][210] = in_1[210] + e1[0][210] %3329;
                                                                                                                                                                                 u[0][211] = in_1[211] + e1[0][211] %3329;
                                                                                                                                                                                 u[0][212] = in_1[212] + e1[0][212] %3329;
                                                                                                                                                                                 u[0][213] = in_1[213] + e1[0][213] %3329;
                                                                                                                                                                                 u[0][214] = in_1[214] + e1[0][214] %3329;
                                                                                                                                                                                 u[0][215] = in_1[215] + e1[0][215] %3329;
                                                                                                                                                                                 u[0][216] = in_1[216] + e1[0][216] %3329;
                                                                                                                                                                                 u[0][217] = in_1[217] + e1[0][217] %3329;
                                                                                                                                                                                 u[0][218] = in_1[218] + e1[0][218] %3329;
                                                                                                                                                                                 u[0][219] = in_1[219] + e1[0][219] %3329;
                                                                                                                                                                                 u[0][220] = in_1[220] + e1[0][220] %3329;
                                                                                                                                                                                 u[0][221] = in_1[221] + e1[0][221] %3329;
                                                                                                                                                                                 u[0][222] = in_1[222] + e1[0][222] %3329;
                                                                                                                                                                                 u[0][223] = in_1[223] + e1[0][223] %3329;
                                                                                                                                                                                 u[0][224] = in_1[224] + e1[0][224] %3329;
                                                                                                                                                                                 u[0][225] = in_1[225] + e1[0][225] %3329;
                                                                                                                                                                                 u[0][226] = in_1[226] + e1[0][226] %3329;
                                                                                                                                                                                 u[0][227] = in_1[227] + e1[0][227] %3329;
                                                                                                                                                                                 u[0][228] = in_1[228] + e1[0][228] %3329;
                                                                                                                                                                                 u[0][229] = in_1[229] + e1[0][229] %3329;
                                                                                                                                                                                 u[0][230] = in_1[230] + e1[0][230] %3329;
                                                                                                                                                                                 u[0][231] = in_1[231] + e1[0][231] %3329;
                                                                                                                                                                                 u[0][232] = in_1[232] + e1[0][232] %3329;
                                                                                                                                                                                 u[0][233] = in_1[233] + e1[0][233] %3329;
                                                                                                                                                                                 u[0][234] = in_1[234] + e1[0][234] %3329;
                                                                                                                                                                                 u[0][235] = in_1[235] + e1[0][235] %3329;
                                                                                                                                                                                 u[0][236] = in_1[236] + e1[0][236] %3329;
                                                                                                                                                                                 u[0][237] = in_1[237] + e1[0][237] %3329;
                                                                                                                                                                                 u[0][238] = in_1[238] + e1[0][238] %3329;
                                                                                                                                                                                 u[0][239] = in_1[239] + e1[0][239] %3329;
                                                                                                                                                                                 u[0][240] = in_1[240] + e1[0][240] %3329;
                                                                                                                                                                                 u[0][241] = in_1[241] + e1[0][241] %3329;
                                                                                                                                                                                 u[0][242] = in_1[242] + e1[0][242] %3329;
                                                                                                                                                                                 u[0][243] = in_1[243] + e1[0][243] %3329;
                                                                                                                                                                                 u[0][244] = in_1[244] + e1[0][244] %3329;
                                                                                                                                                                                 u[0][245] = in_1[245] + e1[0][245] %3329;
                                                                                                                                                                                 u[0][246] = in_1[246] + e1[0][246] %3329;
                                                                                                                                                                                 u[0][247] = in_1[247] + e1[0][247] %3329;
                                                                                                                                                                                 u[0][248] = in_1[248] + e1[0][248] %3329;
                                                                                                                                                                                 u[0][249] = in_1[249] + e1[0][249] %3329;
                                                                                                                                                                                 u[0][250] = in_1[250] + e1[0][250] %3329;
                                                                                                                                                                                 u[0][251] = in_1[251] + e1[0][251] %3329;
                                                                                                                                                                                 u[0][252] = in_1[252] + e1[0][252] %3329;
                                                                                                                                                                                 u[0][253] = in_1[253] + e1[0][253] %3329;
                                                                                                                                                                                 u[0][254] = in_1[254] + e1[0][254] %3329;
                                                                                                                                                                                 u[0][255] = in_1[255] + e1[0][255] %3329;
                                                                                                                                                                                 u[1][0] = in_2[0] + e1[1][0] %3329;
                                                                                                                                                                                 u[1][1] = in_2[1] + e1[1][1] %3329;
                                                                                                                                                                                 u[1][2] = in_2[2] + e1[1][2] %3329;
                                                                                                                                                                                 u[1][3] = in_2[3] + e1[1][3] %3329;
                                                                                                                                                                                 u[1][4] = in_2[4] + e1[1][4] %3329;
                                                                                                                                                                                 u[1][5] = in_2[5] + e1[1][5] %3329;
                                                                                                                                                                                 u[1][6] = in_2[6] + e1[1][6] %3329;
                                                                                                                                                                                 u[1][7] = in_2[7] + e1[1][7] %3329;
                                                                                                                                                                                 u[1][8] = in_2[8] + e1[1][8] %3329;
                                                                                                                                                                                 u[1][9] = in_2[9] + e1[1][9] %3329;
                                                                                                                                                                                 u[1][10] = in_2[10] + e1[1][10] %3329;
                                                                                                                                                                                 u[1][11] = in_2[11] + e1[1][11] %3329;
                                                                                                                                                                                 u[1][12] = in_2[12] + e1[1][12] %3329;
                                                                                                                                                                                 u[1][13] = in_2[13] + e1[1][13] %3329;
                                                                                                                                                                                 u[1][14] = in_2[14] + e1[1][14] %3329;
                                                                                                                                                                                 u[1][15] = in_2[15] + e1[1][15] %3329;
                                                                                                                                                                                 u[1][16] = in_2[16] + e1[1][16] %3329;
                                                                                                                                                                                 u[1][17] = in_2[17] + e1[1][17] %3329;
                                                                                                                                                                                 u[1][18] = in_2[18] + e1[1][18] %3329;
                                                                                                                                                                                 u[1][19] = in_2[19] + e1[1][19] %3329;
                                                                                                                                                                                 u[1][20] = in_2[20] + e1[1][20] %3329;
                                                                                                                                                                                 u[1][21] = in_2[21] + e1[1][21] %3329;
                                                                                                                                                                                 u[1][22] = in_2[22] + e1[1][22] %3329;
                                                                                                                                                                                 u[1][23] = in_2[23] + e1[1][23] %3329;
                                                                                                                                                                                 u[1][24] = in_2[24] + e1[1][24] %3329;
                                                                                                                                                                                 u[1][25] = in_2[25] + e1[1][25] %3329;
                                                                                                                                                                                 u[1][26] = in_2[26] + e1[1][26] %3329;
                                                                                                                                                                                 u[1][27] = in_2[27] + e1[1][27] %3329;
                                                                                                                                                                                 u[1][28] = in_2[28] + e1[1][28] %3329;
                                                                                                                                                                                 u[1][29] = in_2[29] + e1[1][29] %3329;
                                                                                                                                                                                 u[1][30] = in_2[30] + e1[1][30] %3329;
                                                                                                                                                                                 u[1][31] = in_2[31] + e1[1][31] %3329;
                                                                                                                                                                                 u[1][32] = in_2[32] + e1[1][32] %3329;
                                                                                                                                                                                 u[1][33] = in_2[33] + e1[1][33] %3329;
                                                                                                                                                                                 u[1][34] = in_2[34] + e1[1][34] %3329;
                                                                                                                                                                                 u[1][35] = in_2[35] + e1[1][35] %3329;
                                                                                                                                                                                 u[1][36] = in_2[36] + e1[1][36] %3329;
                                                                                                                                                                                 u[1][37] = in_2[37] + e1[1][37] %3329;
                                                                                                                                                                                 u[1][38] = in_2[38] + e1[1][38] %3329;
                                                                                                                                                                                 u[1][39] = in_2[39] + e1[1][39] %3329;
                                                                                                                                                                                 u[1][40] = in_2[40] + e1[1][40] %3329;
                                                                                                                                                                                 u[1][41] = in_2[41] + e1[1][41] %3329;
                                                                                                                                                                                 u[1][42] = in_2[42] + e1[1][42] %3329;
                                                                                                                                                                                 u[1][43] = in_2[43] + e1[1][43] %3329;
                                                                                                                                                                                 u[1][44] = in_2[44] + e1[1][44] %3329;
                                                                                                                                                                                 u[1][45] = in_2[45] + e1[1][45] %3329;
                                                                                                                                                                                 u[1][46] = in_2[46] + e1[1][46] %3329;
                                                                                                                                                                                 u[1][47] = in_2[47] + e1[1][47] %3329;
                                                                                                                                                                                 u[1][48] = in_2[48] + e1[1][48] %3329;
                                                                                                                                                                                 u[1][49] = in_2[49] + e1[1][49] %3329;
                                                                                                                                                                                 u[1][50] = in_2[50] + e1[1][50] %3329;
                                                                                                                                                                                 u[1][51] = in_2[51] + e1[1][51] %3329;
                                                                                                                                                                                 u[1][52] = in_2[52] + e1[1][52] %3329;
                                                                                                                                                                                 u[1][53] = in_2[53] + e1[1][53] %3329;
                                                                                                                                                                                 u[1][54] = in_2[54] + e1[1][54] %3329;
                                                                                                                                                                                 u[1][55] = in_2[55] + e1[1][55] %3329;
                                                                                                                                                                                 u[1][56] = in_2[56] + e1[1][56] %3329;
                                                                                                                                                                                 u[1][57] = in_2[57] + e1[1][57] %3329;
                                                                                                                                                                                 u[1][58] = in_2[58] + e1[1][58] %3329;
                                                                                                                                                                                 u[1][59] = in_2[59] + e1[1][59] %3329;
                                                                                                                                                                                 u[1][60] = in_2[60] + e1[1][60] %3329;
                                                                                                                                                                                 u[1][61] = in_2[61] + e1[1][61] %3329;
                                                                                                                                                                                 u[1][62] = in_2[62] + e1[1][62] %3329;
                                                                                                                                                                                 u[1][63] = in_2[63] + e1[1][63] %3329;
                                                                                                                                                                                 u[1][64] = in_2[64] + e1[1][64] %3329;
                                                                                                                                                                                 u[1][65] = in_2[65] + e1[1][65] %3329;
                                                                                                                                                                                 u[1][66] = in_2[66] + e1[1][66] %3329;
                                                                                                                                                                                 u[1][67] = in_2[67] + e1[1][67] %3329;
                                                                                                                                                                                 u[1][68] = in_2[68] + e1[1][68] %3329;
                                                                                                                                                                                 u[1][69] = in_2[69] + e1[1][69] %3329;
                                                                                                                                                                                 u[1][70] = in_2[70] + e1[1][70] %3329;
                                                                                                                                                                                 u[1][71] = in_2[71] + e1[1][71] %3329;
                                                                                                                                                                                 u[1][72] = in_2[72] + e1[1][72] %3329;
                                                                                                                                                                                 u[1][73] = in_2[73] + e1[1][73] %3329;
                                                                                                                                                                                 u[1][74] = in_2[74] + e1[1][74] %3329;
                                                                                                                                                                                 u[1][75] = in_2[75] + e1[1][75] %3329;
                                                                                                                                                                                 u[1][76] = in_2[76] + e1[1][76] %3329;
                                                                                                                                                                                 u[1][77] = in_2[77] + e1[1][77] %3329;
                                                                                                                                                                                 u[1][78] = in_2[78] + e1[1][78] %3329;
                                                                                                                                                                                 u[1][79] = in_2[79] + e1[1][79] %3329;
                                                                                                                                                                                 u[1][80] = in_2[80] + e1[1][80] %3329;
                                                                                                                                                                                 u[1][81] = in_2[81] + e1[1][81] %3329;
                                                                                                                                                                                 u[1][82] = in_2[82] + e1[1][82] %3329;
                                                                                                                                                                                 u[1][83] = in_2[83] + e1[1][83] %3329;
                                                                                                                                                                                 u[1][84] = in_2[84] + e1[1][84] %3329;
                                                                                                                                                                                 u[1][85] = in_2[85] + e1[1][85] %3329;
                                                                                                                                                                                 u[1][86] = in_2[86] + e1[1][86] %3329;
                                                                                                                                                                                 u[1][87] = in_2[87] + e1[1][87] %3329;
                                                                                                                                                                                 u[1][88] = in_2[88] + e1[1][88] %3329;
                                                                                                                                                                                 u[1][89] = in_2[89] + e1[1][89] %3329;
                                                                                                                                                                                 u[1][90] = in_2[90] + e1[1][90] %3329;
                                                                                                                                                                                 u[1][91] = in_2[91] + e1[1][91] %3329;
                                                                                                                                                                                 u[1][92] = in_2[92] + e1[1][92] %3329;
                                                                                                                                                                                 u[1][93] = in_2[93] + e1[1][93] %3329;
                                                                                                                                                                                 u[1][94] = in_2[94] + e1[1][94] %3329;
                                                                                                                                                                                 u[1][95] = in_2[95] + e1[1][95] %3329;
                                                                                                                                                                                 u[1][96] = in_2[96] + e1[1][96] %3329;
                                                                                                                                                                                 u[1][97] = in_2[97] + e1[1][97] %3329;
                                                                                                                                                                                 u[1][98] = in_2[98] + e1[1][98] %3329;
                                                                                                                                                                                 u[1][99] = in_2[99] + e1[1][99] %3329;
                                                                                                                                                                                 u[1][100] = in_2[100] + e1[1][100] %3329;
                                                                                                                                                                                 u[1][101] = in_2[101] + e1[1][101] %3329;
                                                                                                                                                                                 u[1][102] = in_2[102] + e1[1][102] %3329;
                                                                                                                                                                                 u[1][103] = in_2[103] + e1[1][103] %3329;
                                                                                                                                                                                 u[1][104] = in_2[104] + e1[1][104] %3329;
                                                                                                                                                                                 u[1][105] = in_2[105] + e1[1][105] %3329;
                                                                                                                                                                                 u[1][106] = in_2[106] + e1[1][106] %3329;
                                                                                                                                                                                 u[1][107] = in_2[107] + e1[1][107] %3329;
                                                                                                                                                                                 u[1][108] = in_2[108] + e1[1][108] %3329;
                                                                                                                                                                                 u[1][109] = in_2[109] + e1[1][109] %3329;
                                                                                                                                                                                 u[1][110] = in_2[110] + e1[1][110] %3329;
                                                                                                                                                                                 u[1][111] = in_2[111] + e1[1][111] %3329;
                                                                                                                                                                                 u[1][112] = in_2[112] + e1[1][112] %3329;
                                                                                                                                                                                 u[1][113] = in_2[113] + e1[1][113] %3329;
                                                                                                                                                                                 u[1][114] = in_2[114] + e1[1][114] %3329;
                                                                                                                                                                                 u[1][115] = in_2[115] + e1[1][115] %3329;
                                                                                                                                                                                 u[1][116] = in_2[116] + e1[1][116] %3329;
                                                                                                                                                                                 u[1][117] = in_2[117] + e1[1][117] %3329;
                                                                                                                                                                                 u[1][118] = in_2[118] + e1[1][118] %3329;
                                                                                                                                                                                 u[1][119] = in_2[119] + e1[1][119] %3329;
                                                                                                                                                                                 u[1][120] = in_2[120] + e1[1][120] %3329;
                                                                                                                                                                                 u[1][121] = in_2[121] + e1[1][121] %3329;
                                                                                                                                                                                 u[1][122] = in_2[122] + e1[1][122] %3329;
                                                                                                                                                                                 u[1][123] = in_2[123] + e1[1][123] %3329;
                                                                                                                                                                                 u[1][124] = in_2[124] + e1[1][124] %3329;
                                                                                                                                                                                 u[1][125] = in_2[125] + e1[1][125] %3329;
                                                                                                                                                                                 u[1][126] = in_2[126] + e1[1][126] %3329;
                                                                                                                                                                                 u[1][127] = in_2[127] + e1[1][127] %3329;
                                                                                                                                                                                 u[1][128] = in_2[128] + e1[1][128] %3329;
                                                                                                                                                                                 u[1][129] = in_2[129] + e1[1][129] %3329;
                                                                                                                                                                                 u[1][130] = in_2[130] + e1[1][130] %3329;
                                                                                                                                                                                 u[1][131] = in_2[131] + e1[1][131] %3329;
                                                                                                                                                                                 u[1][132] = in_2[132] + e1[1][132] %3329;
                                                                                                                                                                                 u[1][133] = in_2[133] + e1[1][133] %3329;
                                                                                                                                                                                 u[1][134] = in_2[134] + e1[1][134] %3329;
                                                                                                                                                                                 u[1][135] = in_2[135] + e1[1][135] %3329;
                                                                                                                                                                                 u[1][136] = in_2[136] + e1[1][136] %3329;
                                                                                                                                                                                 u[1][137] = in_2[137] + e1[1][137] %3329;
                                                                                                                                                                                 u[1][138] = in_2[138] + e1[1][138] %3329;
                                                                                                                                                                                 u[1][139] = in_2[139] + e1[1][139] %3329;
                                                                                                                                                                                 u[1][140] = in_2[140] + e1[1][140] %3329;
                                                                                                                                                                                 u[1][141] = in_2[141] + e1[1][141] %3329;
                                                                                                                                                                                 u[1][142] = in_2[142] + e1[1][142] %3329;
                                                                                                                                                                                 u[1][143] = in_2[143] + e1[1][143] %3329;
                                                                                                                                                                                 u[1][144] = in_2[144] + e1[1][144] %3329;
                                                                                                                                                                                 u[1][145] = in_2[145] + e1[1][145] %3329;
                                                                                                                                                                                 u[1][146] = in_2[146] + e1[1][146] %3329;
                                                                                                                                                                                 u[1][147] = in_2[147] + e1[1][147] %3329;
                                                                                                                                                                                 u[1][148] = in_2[148] + e1[1][148] %3329;
                                                                                                                                                                                 u[1][149] = in_2[149] + e1[1][149] %3329;
                                                                                                                                                                                 u[1][150] = in_2[150] + e1[1][150] %3329;
                                                                                                                                                                                 u[1][151] = in_2[151] + e1[1][151] %3329;
                                                                                                                                                                                 u[1][152] = in_2[152] + e1[1][152] %3329;
                                                                                                                                                                                 u[1][153] = in_2[153] + e1[1][153] %3329;
                                                                                                                                                                                 u[1][154] = in_2[154] + e1[1][154] %3329;
                                                                                                                                                                                 u[1][155] = in_2[155] + e1[1][155] %3329;
                                                                                                                                                                                 u[1][156] = in_2[156] + e1[1][156] %3329;
                                                                                                                                                                                 u[1][157] = in_2[157] + e1[1][157] %3329;
                                                                                                                                                                                 u[1][158] = in_2[158] + e1[1][158] %3329;
                                                                                                                                                                                 u[1][159] = in_2[159] + e1[1][159] %3329;
                                                                                                                                                                                 u[1][160] = in_2[160] + e1[1][160] %3329;
                                                                                                                                                                                 u[1][161] = in_2[161] + e1[1][161] %3329;
                                                                                                                                                                                 u[1][162] = in_2[162] + e1[1][162] %3329;
                                                                                                                                                                                 u[1][163] = in_2[163] + e1[1][163] %3329;
                                                                                                                                                                                 u[1][164] = in_2[164] + e1[1][164] %3329;
                                                                                                                                                                                 u[1][165] = in_2[165] + e1[1][165] %3329;
                                                                                                                                                                                 u[1][166] = in_2[166] + e1[1][166] %3329;
                                                                                                                                                                                 u[1][167] = in_2[167] + e1[1][167] %3329;
                                                                                                                                                                                 u[1][168] = in_2[168] + e1[1][168] %3329;
                                                                                                                                                                                 u[1][169] = in_2[169] + e1[1][169] %3329;
                                                                                                                                                                                 u[1][170] = in_2[170] + e1[1][170] %3329;
                                                                                                                                                                                 u[1][171] = in_2[171] + e1[1][171] %3329;
                                                                                                                                                                                 u[1][172] = in_2[172] + e1[1][172] %3329;
                                                                                                                                                                                 u[1][173] = in_2[173] + e1[1][173] %3329;
                                                                                                                                                                                 u[1][174] = in_2[174] + e1[1][174] %3329;
                                                                                                                                                                                 u[1][175] = in_2[175] + e1[1][175] %3329;
                                                                                                                                                                                 u[1][176] = in_2[176] + e1[1][176] %3329;
                                                                                                                                                                                 u[1][177] = in_2[177] + e1[1][177] %3329;
                                                                                                                                                                                 u[1][178] = in_2[178] + e1[1][178] %3329;
                                                                                                                                                                                 u[1][179] = in_2[179] + e1[1][179] %3329;
                                                                                                                                                                                 u[1][180] = in_2[180] + e1[1][180] %3329;
                                                                                                                                                                                 u[1][181] = in_2[181] + e1[1][181] %3329;
                                                                                                                                                                                 u[1][182] = in_2[182] + e1[1][182] %3329;
                                                                                                                                                                                 u[1][183] = in_2[183] + e1[1][183] %3329;
                                                                                                                                                                                 u[1][184] = in_2[184] + e1[1][184] %3329;
                                                                                                                                                                                 u[1][185] = in_2[185] + e1[1][185] %3329;
                                                                                                                                                                                 u[1][186] = in_2[186] + e1[1][186] %3329;
                                                                                                                                                                                 u[1][187] = in_2[187] + e1[1][187] %3329;
                                                                                                                                                                                 u[1][188] = in_2[188] + e1[1][188] %3329;
                                                                                                                                                                                 u[1][189] = in_2[189] + e1[1][189] %3329;
                                                                                                                                                                                 u[1][190] = in_2[190] + e1[1][190] %3329;
                                                                                                                                                                                 u[1][191] = in_2[191] + e1[1][191] %3329;
                                                                                                                                                                                 u[1][192] = in_2[192] + e1[1][192] %3329;
                                                                                                                                                                                 u[1][193] = in_2[193] + e1[1][193] %3329;
                                                                                                                                                                                 u[1][194] = in_2[194] + e1[1][194] %3329;
                                                                                                                                                                                 u[1][195] = in_2[195] + e1[1][195] %3329;
                                                                                                                                                                                 u[1][196] = in_2[196] + e1[1][196] %3329;
                                                                                                                                                                                 u[1][197] = in_2[197] + e1[1][197] %3329;
                                                                                                                                                                                 u[1][198] = in_2[198] + e1[1][198] %3329;
                                                                                                                                                                                 u[1][199] = in_2[199] + e1[1][199] %3329;
                                                                                                                                                                                 u[1][200] = in_2[200] + e1[1][200] %3329;
                                                                                                                                                                                 u[1][201] = in_2[201] + e1[1][201] %3329;
                                                                                                                                                                                 u[1][202] = in_2[202] + e1[1][202] %3329;
                                                                                                                                                                                 u[1][203] = in_2[203] + e1[1][203] %3329;
                                                                                                                                                                                 u[1][204] = in_2[204] + e1[1][204] %3329;
                                                                                                                                                                                 u[1][205] = in_2[205] + e1[1][205] %3329;
                                                                                                                                                                                 u[1][206] = in_2[206] + e1[1][206] %3329;
                                                                                                                                                                                 u[1][207] = in_2[207] + e1[1][207] %3329;
                                                                                                                                                                                 u[1][208] = in_2[208] + e1[1][208] %3329;
                                                                                                                                                                                 u[1][209] = in_2[209] + e1[1][209] %3329;
                                                                                                                                                                                 u[1][210] = in_2[210] + e1[1][210] %3329;
                                                                                                                                                                                 u[1][211] = in_2[211] + e1[1][211] %3329;
                                                                                                                                                                                 u[1][212] = in_2[212] + e1[1][212] %3329;
                                                                                                                                                                                 u[1][213] = in_2[213] + e1[1][213] %3329;
                                                                                                                                                                                 u[1][214] = in_2[214] + e1[1][214] %3329;
                                                                                                                                                                                 u[1][215] = in_2[215] + e1[1][215] %3329;
                                                                                                                                                                                 u[1][216] = in_2[216] + e1[1][216] %3329;
                                                                                                                                                                                 u[1][217] = in_2[217] + e1[1][217] %3329;
                                                                                                                                                                                 u[1][218] = in_2[218] + e1[1][218] %3329;
                                                                                                                                                                                 u[1][219] = in_2[219] + e1[1][219] %3329;
                                                                                                                                                                                 u[1][220] = in_2[220] + e1[1][220] %3329;
                                                                                                                                                                                 u[1][221] = in_2[221] + e1[1][221] %3329;
                                                                                                                                                                                 u[1][222] = in_2[222] + e1[1][222] %3329;
                                                                                                                                                                                 u[1][223] = in_2[223] + e1[1][223] %3329;
                                                                                                                                                                                 u[1][224] = in_2[224] + e1[1][224] %3329;
                                                                                                                                                                                 u[1][225] = in_2[225] + e1[1][225] %3329;
                                                                                                                                                                                 u[1][226] = in_2[226] + e1[1][226] %3329;
                                                                                                                                                                                 u[1][227] = in_2[227] + e1[1][227] %3329;
                                                                                                                                                                                 u[1][228] = in_2[228] + e1[1][228] %3329;
                                                                                                                                                                                 u[1][229] = in_2[229] + e1[1][229] %3329;
                                                                                                                                                                                 u[1][230] = in_2[230] + e1[1][230] %3329;
                                                                                                                                                                                 u[1][231] = in_2[231] + e1[1][231] %3329;
                                                                                                                                                                                 u[1][232] = in_2[232] + e1[1][232] %3329;
                                                                                                                                                                                 u[1][233] = in_2[233] + e1[1][233] %3329;
                                                                                                                                                                                 u[1][234] = in_2[234] + e1[1][234] %3329;
                                                                                                                                                                                 u[1][235] = in_2[235] + e1[1][235] %3329;
                                                                                                                                                                                 u[1][236] = in_2[236] + e1[1][236] %3329;
                                                                                                                                                                                 u[1][237] = in_2[237] + e1[1][237] %3329;
                                                                                                                                                                                 u[1][238] = in_2[238] + e1[1][238] %3329;
                                                                                                                                                                                 u[1][239] = in_2[239] + e1[1][239] %3329;
                                                                                                                                                                                 u[1][240] = in_2[240] + e1[1][240] %3329;
                                                                                                                                                                                 u[1][241] = in_2[241] + e1[1][241] %3329;
                                                                                                                                                                                 u[1][242] = in_2[242] + e1[1][242] %3329;
                                                                                                                                                                                 u[1][243] = in_2[243] + e1[1][243] %3329;
                                                                                                                                                                                 u[1][244] = in_2[244] + e1[1][244] %3329;
                                                                                                                                                                                 u[1][245] = in_2[245] + e1[1][245] %3329;
                                                                                                                                                                                 u[1][246] = in_2[246] + e1[1][246] %3329;
                                                                                                                                                                                 u[1][247] = in_2[247] + e1[1][247] %3329;
                                                                                                                                                                                 u[1][248] = in_2[248] + e1[1][248] %3329;
                                                                                                                                                                                 u[1][249] = in_2[249] + e1[1][249] %3329;
                                                                                                                                                                                 u[1][250] = in_2[250] + e1[1][250] %3329;
                                                                                                                                                                                 u[1][251] = in_2[251] + e1[1][251] %3329;
                                                                                                                                                                                 u[1][252] = in_2[252] + e1[1][252] %3329;
                                                                                                                                                                                 u[1][253] = in_2[253] + e1[1][253] %3329;
                                                                                                                                                                                 u[1][254] = in_2[254] + e1[1][254] %3329;
                                                                                                                                                                                 u[1][255] = in_2[255] + e1[1][255] %3329;
                                                                                                                                                                                 u[2][0] = in_3[0] + e1[2][0] %3329;
                                                                                                                                                                                 u[2][1] = in_3[1] + e1[2][1] %3329;
                                                                                                                                                                                 u[2][2] = in_3[2] + e1[2][2] %3329;
                                                                                                                                                                                 u[2][3] = in_3[3] + e1[2][3] %3329;
                                                                                                                                                                                 u[2][4] = in_3[4] + e1[2][4] %3329;
                                                                                                                                                                                 u[2][5] = in_3[5] + e1[2][5] %3329;
                                                                                                                                                                                 u[2][6] = in_3[6] + e1[2][6] %3329;
                                                                                                                                                                                 u[2][7] = in_3[7] + e1[2][7] %3329;
                                                                                                                                                                                 u[2][8] = in_3[8] + e1[2][8] %3329;
                                                                                                                                                                                 u[2][9] = in_3[9] + e1[2][9] %3329;
                                                                                                                                                                                 u[2][10] = in_3[10] + e1[2][10] %3329;
                                                                                                                                                                                 u[2][11] = in_3[11] + e1[2][11] %3329;
                                                                                                                                                                                 u[2][12] = in_3[12] + e1[2][12] %3329;
                                                                                                                                                                                 u[2][13] = in_3[13] + e1[2][13] %3329;
                                                                                                                                                                                 u[2][14] = in_3[14] + e1[2][14] %3329;
                                                                                                                                                                                 u[2][15] = in_3[15] + e1[2][15] %3329;
                                                                                                                                                                                 u[2][16] = in_3[16] + e1[2][16] %3329;
                                                                                                                                                                                 u[2][17] = in_3[17] + e1[2][17] %3329;
                                                                                                                                                                                 u[2][18] = in_3[18] + e1[2][18] %3329;
                                                                                                                                                                                 u[2][19] = in_3[19] + e1[2][19] %3329;
                                                                                                                                                                                 u[2][20] = in_3[20] + e1[2][20] %3329;
                                                                                                                                                                                 u[2][21] = in_3[21] + e1[2][21] %3329;
                                                                                                                                                                                 u[2][22] = in_3[22] + e1[2][22] %3329;
                                                                                                                                                                                 u[2][23] = in_3[23] + e1[2][23] %3329;
                                                                                                                                                                                 u[2][24] = in_3[24] + e1[2][24] %3329;
                                                                                                                                                                                 u[2][25] = in_3[25] + e1[2][25] %3329;
                                                                                                                                                                                 u[2][26] = in_3[26] + e1[2][26] %3329;
                                                                                                                                                                                 u[2][27] = in_3[27] + e1[2][27] %3329;
                                                                                                                                                                                 u[2][28] = in_3[28] + e1[2][28] %3329;
                                                                                                                                                                                 u[2][29] = in_3[29] + e1[2][29] %3329;
                                                                                                                                                                                 u[2][30] = in_3[30] + e1[2][30] %3329;
                                                                                                                                                                                 u[2][31] = in_3[31] + e1[2][31] %3329;
                                                                                                                                                                                 u[2][32] = in_3[32] + e1[2][32] %3329;
                                                                                                                                                                                 u[2][33] = in_3[33] + e1[2][33] %3329;
                                                                                                                                                                                 u[2][34] = in_3[34] + e1[2][34] %3329;
                                                                                                                                                                                 u[2][35] = in_3[35] + e1[2][35] %3329;
                                                                                                                                                                                 u[2][36] = in_3[36] + e1[2][36] %3329;
                                                                                                                                                                                 u[2][37] = in_3[37] + e1[2][37] %3329;
                                                                                                                                                                                 u[2][38] = in_3[38] + e1[2][38] %3329;
                                                                                                                                                                                 u[2][39] = in_3[39] + e1[2][39] %3329;
                                                                                                                                                                                 u[2][40] = in_3[40] + e1[2][40] %3329;
                                                                                                                                                                                 u[2][41] = in_3[41] + e1[2][41] %3329;
                                                                                                                                                                                 u[2][42] = in_3[42] + e1[2][42] %3329;
                                                                                                                                                                                 u[2][43] = in_3[43] + e1[2][43] %3329;
                                                                                                                                                                                 u[2][44] = in_3[44] + e1[2][44] %3329;
                                                                                                                                                                                 u[2][45] = in_3[45] + e1[2][45] %3329;
                                                                                                                                                                                 u[2][46] = in_3[46] + e1[2][46] %3329;
                                                                                                                                                                                 u[2][47] = in_3[47] + e1[2][47] %3329;
                                                                                                                                                                                 u[2][48] = in_3[48] + e1[2][48] %3329;
                                                                                                                                                                                 u[2][49] = in_3[49] + e1[2][49] %3329;
                                                                                                                                                                                 u[2][50] = in_3[50] + e1[2][50] %3329;
                                                                                                                                                                                 u[2][51] = in_3[51] + e1[2][51] %3329;
                                                                                                                                                                                 u[2][52] = in_3[52] + e1[2][52] %3329;
                                                                                                                                                                                 u[2][53] = in_3[53] + e1[2][53] %3329;
                                                                                                                                                                                 u[2][54] = in_3[54] + e1[2][54] %3329;
                                                                                                                                                                                 u[2][55] = in_3[55] + e1[2][55] %3329;
                                                                                                                                                                                 u[2][56] = in_3[56] + e1[2][56] %3329;
                                                                                                                                                                                 u[2][57] = in_3[57] + e1[2][57] %3329;
                                                                                                                                                                                 u[2][58] = in_3[58] + e1[2][58] %3329;
                                                                                                                                                                                 u[2][59] = in_3[59] + e1[2][59] %3329;
                                                                                                                                                                                 u[2][60] = in_3[60] + e1[2][60] %3329;
                                                                                                                                                                                 u[2][61] = in_3[61] + e1[2][61] %3329;
                                                                                                                                                                                 u[2][62] = in_3[62] + e1[2][62] %3329;
                                                                                                                                                                                 u[2][63] = in_3[63] + e1[2][63] %3329;
                                                                                                                                                                                 u[2][64] = in_3[64] + e1[2][64] %3329;
                                                                                                                                                                                 u[2][65] = in_3[65] + e1[2][65] %3329;
                                                                                                                                                                                 u[2][66] = in_3[66] + e1[2][66] %3329;
                                                                                                                                                                                 u[2][67] = in_3[67] + e1[2][67] %3329;
                                                                                                                                                                                 u[2][68] = in_3[68] + e1[2][68] %3329;
                                                                                                                                                                                 u[2][69] = in_3[69] + e1[2][69] %3329;
                                                                                                                                                                                 u[2][70] = in_3[70] + e1[2][70] %3329;
                                                                                                                                                                                 u[2][71] = in_3[71] + e1[2][71] %3329;
                                                                                                                                                                                 u[2][72] = in_3[72] + e1[2][72] %3329;
                                                                                                                                                                                 u[2][73] = in_3[73] + e1[2][73] %3329;
                                                                                                                                                                                 u[2][74] = in_3[74] + e1[2][74] %3329;
                                                                                                                                                                                 u[2][75] = in_3[75] + e1[2][75] %3329;
                                                                                                                                                                                 u[2][76] = in_3[76] + e1[2][76] %3329;
                                                                                                                                                                                 u[2][77] = in_3[77] + e1[2][77] %3329;
                                                                                                                                                                                 u[2][78] = in_3[78] + e1[2][78] %3329;
                                                                                                                                                                                 u[2][79] = in_3[79] + e1[2][79] %3329;
                                                                                                                                                                                 u[2][80] = in_3[80] + e1[2][80] %3329;
                                                                                                                                                                                 u[2][81] = in_3[81] + e1[2][81] %3329;
                                                                                                                                                                                 u[2][82] = in_3[82] + e1[2][82] %3329;
                                                                                                                                                                                 u[2][83] = in_3[83] + e1[2][83] %3329;
                                                                                                                                                                                 u[2][84] = in_3[84] + e1[2][84] %3329;
                                                                                                                                                                                 u[2][85] = in_3[85] + e1[2][85] %3329;
                                                                                                                                                                                 u[2][86] = in_3[86] + e1[2][86] %3329;
                                                                                                                                                                                 u[2][87] = in_3[87] + e1[2][87] %3329;
                                                                                                                                                                                 u[2][88] = in_3[88] + e1[2][88] %3329;
                                                                                                                                                                                 u[2][89] = in_3[89] + e1[2][89] %3329;
                                                                                                                                                                                 u[2][90] = in_3[90] + e1[2][90] %3329;
                                                                                                                                                                                 u[2][91] = in_3[91] + e1[2][91] %3329;
                                                                                                                                                                                 u[2][92] = in_3[92] + e1[2][92] %3329;
                                                                                                                                                                                 u[2][93] = in_3[93] + e1[2][93] %3329;
                                                                                                                                                                                 u[2][94] = in_3[94] + e1[2][94] %3329;
                                                                                                                                                                                 u[2][95] = in_3[95] + e1[2][95] %3329;
                                                                                                                                                                                 u[2][96] = in_3[96] + e1[2][96] %3329;
                                                                                                                                                                                 u[2][97] = in_3[97] + e1[2][97] %3329;
                                                                                                                                                                                 u[2][98] = in_3[98] + e1[2][98] %3329;
                                                                                                                                                                                 u[2][99] = in_3[99] + e1[2][99] %3329;
                                                                                                                                                                                 u[2][100] = in_3[100] + e1[2][100] %3329;
                                                                                                                                                                                 u[2][101] = in_3[101] + e1[2][101] %3329;
                                                                                                                                                                                 u[2][102] = in_3[102] + e1[2][102] %3329;
                                                                                                                                                                                 u[2][103] = in_3[103] + e1[2][103] %3329;
                                                                                                                                                                                 u[2][104] = in_3[104] + e1[2][104] %3329;
                                                                                                                                                                                 u[2][105] = in_3[105] + e1[2][105] %3329;
                                                                                                                                                                                 u[2][106] = in_3[106] + e1[2][106] %3329;
                                                                                                                                                                                 u[2][107] = in_3[107] + e1[2][107] %3329;
                                                                                                                                                                                 u[2][108] = in_3[108] + e1[2][108] %3329;
                                                                                                                                                                                 u[2][109] = in_3[109] + e1[2][109] %3329;
                                                                                                                                                                                 u[2][110] = in_3[110] + e1[2][110] %3329;
                                                                                                                                                                                 u[2][111] = in_3[111] + e1[2][111] %3329;
                                                                                                                                                                                 u[2][112] = in_3[112] + e1[2][112] %3329;
                                                                                                                                                                                 u[2][113] = in_3[113] + e1[2][113] %3329;
                                                                                                                                                                                 u[2][114] = in_3[114] + e1[2][114] %3329;
                                                                                                                                                                                 u[2][115] = in_3[115] + e1[2][115] %3329;
                                                                                                                                                                                 u[2][116] = in_3[116] + e1[2][116] %3329;
                                                                                                                                                                                 u[2][117] = in_3[117] + e1[2][117] %3329;
                                                                                                                                                                                 u[2][118] = in_3[118] + e1[2][118] %3329;
                                                                                                                                                                                 u[2][119] = in_3[119] + e1[2][119] %3329;
                                                                                                                                                                                 u[2][120] = in_3[120] + e1[2][120] %3329;
                                                                                                                                                                                 u[2][121] = in_3[121] + e1[2][121] %3329;
                                                                                                                                                                                 u[2][122] = in_3[122] + e1[2][122] %3329;
                                                                                                                                                                                 u[2][123] = in_3[123] + e1[2][123] %3329;
                                                                                                                                                                                 u[2][124] = in_3[124] + e1[2][124] %3329;
                                                                                                                                                                                 u[2][125] = in_3[125] + e1[2][125] %3329;
                                                                                                                                                                                 u[2][126] = in_3[126] + e1[2][126] %3329;
                                                                                                                                                                                 u[2][127] = in_3[127] + e1[2][127] %3329;
                                                                                                                                                                                 u[2][128] = in_3[128] + e1[2][128] %3329;
                                                                                                                                                                                 u[2][129] = in_3[129] + e1[2][129] %3329;
                                                                                                                                                                                 u[2][130] = in_3[130] + e1[2][130] %3329;
                                                                                                                                                                                 u[2][131] = in_3[131] + e1[2][131] %3329;
                                                                                                                                                                                 u[2][132] = in_3[132] + e1[2][132] %3329;
                                                                                                                                                                                 u[2][133] = in_3[133] + e1[2][133] %3329;
                                                                                                                                                                                 u[2][134] = in_3[134] + e1[2][134] %3329;
                                                                                                                                                                                 u[2][135] = in_3[135] + e1[2][135] %3329;
                                                                                                                                                                                 u[2][136] = in_3[136] + e1[2][136] %3329;
                                                                                                                                                                                 u[2][137] = in_3[137] + e1[2][137] %3329;
                                                                                                                                                                                 u[2][138] = in_3[138] + e1[2][138] %3329;
                                                                                                                                                                                 u[2][139] = in_3[139] + e1[2][139] %3329;
                                                                                                                                                                                 u[2][140] = in_3[140] + e1[2][140] %3329;
                                                                                                                                                                                 u[2][141] = in_3[141] + e1[2][141] %3329;
                                                                                                                                                                                 u[2][142] = in_3[142] + e1[2][142] %3329;
                                                                                                                                                                                 u[2][143] = in_3[143] + e1[2][143] %3329;
                                                                                                                                                                                 u[2][144] = in_3[144] + e1[2][144] %3329;
                                                                                                                                                                                 u[2][145] = in_3[145] + e1[2][145] %3329;
                                                                                                                                                                                 u[2][146] = in_3[146] + e1[2][146] %3329;
                                                                                                                                                                                 u[2][147] = in_3[147] + e1[2][147] %3329;
                                                                                                                                                                                 u[2][148] = in_3[148] + e1[2][148] %3329;
                                                                                                                                                                                 u[2][149] = in_3[149] + e1[2][149] %3329;
                                                                                                                                                                                 u[2][150] = in_3[150] + e1[2][150] %3329;
                                                                                                                                                                                 u[2][151] = in_3[151] + e1[2][151] %3329;
                                                                                                                                                                                 u[2][152] = in_3[152] + e1[2][152] %3329;
                                                                                                                                                                                 u[2][153] = in_3[153] + e1[2][153] %3329;
                                                                                                                                                                                 u[2][154] = in_3[154] + e1[2][154] %3329;
                                                                                                                                                                                 u[2][155] = in_3[155] + e1[2][155] %3329;
                                                                                                                                                                                 u[2][156] = in_3[156] + e1[2][156] %3329;
                                                                                                                                                                                 u[2][157] = in_3[157] + e1[2][157] %3329;
                                                                                                                                                                                 u[2][158] = in_3[158] + e1[2][158] %3329;
                                                                                                                                                                                 u[2][159] = in_3[159] + e1[2][159] %3329;
                                                                                                                                                                                 u[2][160] = in_3[160] + e1[2][160] %3329;
                                                                                                                                                                                 u[2][161] = in_3[161] + e1[2][161] %3329;
                                                                                                                                                                                 u[2][162] = in_3[162] + e1[2][162] %3329;
                                                                                                                                                                                 u[2][163] = in_3[163] + e1[2][163] %3329;
                                                                                                                                                                                 u[2][164] = in_3[164] + e1[2][164] %3329;
                                                                                                                                                                                 u[2][165] = in_3[165] + e1[2][165] %3329;
                                                                                                                                                                                 u[2][166] = in_3[166] + e1[2][166] %3329;
                                                                                                                                                                                 u[2][167] = in_3[167] + e1[2][167] %3329;
                                                                                                                                                                                 u[2][168] = in_3[168] + e1[2][168] %3329;
                                                                                                                                                                                 u[2][169] = in_3[169] + e1[2][169] %3329;
                                                                                                                                                                                 u[2][170] = in_3[170] + e1[2][170] %3329;
                                                                                                                                                                                 u[2][171] = in_3[171] + e1[2][171] %3329;
                                                                                                                                                                                 u[2][172] = in_3[172] + e1[2][172] %3329;
                                                                                                                                                                                 u[2][173] = in_3[173] + e1[2][173] %3329;
                                                                                                                                                                                 u[2][174] = in_3[174] + e1[2][174] %3329;
                                                                                                                                                                                 u[2][175] = in_3[175] + e1[2][175] %3329;
                                                                                                                                                                                 u[2][176] = in_3[176] + e1[2][176] %3329;
                                                                                                                                                                                 u[2][177] = in_3[177] + e1[2][177] %3329;
                                                                                                                                                                                 u[2][178] = in_3[178] + e1[2][178] %3329;
                                                                                                                                                                                 u[2][179] = in_3[179] + e1[2][179] %3329;
                                                                                                                                                                                 u[2][180] = in_3[180] + e1[2][180] %3329;
                                                                                                                                                                                 u[2][181] = in_3[181] + e1[2][181] %3329;
                                                                                                                                                                                 u[2][182] = in_3[182] + e1[2][182] %3329;
                                                                                                                                                                                 u[2][183] = in_3[183] + e1[2][183] %3329;
                                                                                                                                                                                 u[2][184] = in_3[184] + e1[2][184] %3329;
                                                                                                                                                                                 u[2][185] = in_3[185] + e1[2][185] %3329;
                                                                                                                                                                                 u[2][186] = in_3[186] + e1[2][186] %3329;
                                                                                                                                                                                 u[2][187] = in_3[187] + e1[2][187] %3329;
                                                                                                                                                                                 u[2][188] = in_3[188] + e1[2][188] %3329;
                                                                                                                                                                                 u[2][189] = in_3[189] + e1[2][189] %3329;
                                                                                                                                                                                 u[2][190] = in_3[190] + e1[2][190] %3329;
                                                                                                                                                                                 u[2][191] = in_3[191] + e1[2][191] %3329;
                                                                                                                                                                                 u[2][192] = in_3[192] + e1[2][192] %3329;
                                                                                                                                                                                 u[2][193] = in_3[193] + e1[2][193] %3329;
                                                                                                                                                                                 u[2][194] = in_3[194] + e1[2][194] %3329;
                                                                                                                                                                                 u[2][195] = in_3[195] + e1[2][195] %3329;
                                                                                                                                                                                 u[2][196] = in_3[196] + e1[2][196] %3329;
                                                                                                                                                                                 u[2][197] = in_3[197] + e1[2][197] %3329;
                                                                                                                                                                                 u[2][198] = in_3[198] + e1[2][198] %3329;
                                                                                                                                                                                 u[2][199] = in_3[199] + e1[2][199] %3329;
                                                                                                                                                                                 u[2][200] = in_3[200] + e1[2][200] %3329;
                                                                                                                                                                                 u[2][201] = in_3[201] + e1[2][201] %3329;
                                                                                                                                                                                 u[2][202] = in_3[202] + e1[2][202] %3329;
                                                                                                                                                                                 u[2][203] = in_3[203] + e1[2][203] %3329;
                                                                                                                                                                                 u[2][204] = in_3[204] + e1[2][204] %3329;
                                                                                                                                                                                 u[2][205] = in_3[205] + e1[2][205] %3329;
                                                                                                                                                                                 u[2][206] = in_3[206] + e1[2][206] %3329;
                                                                                                                                                                                 u[2][207] = in_3[207] + e1[2][207] %3329;
                                                                                                                                                                                 u[2][208] = in_3[208] + e1[2][208] %3329;
                                                                                                                                                                                 u[2][209] = in_3[209] + e1[2][209] %3329;
                                                                                                                                                                                 u[2][210] = in_3[210] + e1[2][210] %3329;
                                                                                                                                                                                 u[2][211] = in_3[211] + e1[2][211] %3329;
                                                                                                                                                                                 u[2][212] = in_3[212] + e1[2][212] %3329;
                                                                                                                                                                                 u[2][213] = in_3[213] + e1[2][213] %3329;
                                                                                                                                                                                 u[2][214] = in_3[214] + e1[2][214] %3329;
                                                                                                                                                                                 u[2][215] = in_3[215] + e1[2][215] %3329;
                                                                                                                                                                                 u[2][216] = in_3[216] + e1[2][216] %3329;
                                                                                                                                                                                 u[2][217] = in_3[217] + e1[2][217] %3329;
                                                                                                                                                                                 u[2][218] = in_3[218] + e1[2][218] %3329;
                                                                                                                                                                                 u[2][219] = in_3[219] + e1[2][219] %3329;
                                                                                                                                                                                 u[2][220] = in_3[220] + e1[2][220] %3329;
                                                                                                                                                                                 u[2][221] = in_3[221] + e1[2][221] %3329;
                                                                                                                                                                                 u[2][222] = in_3[222] + e1[2][222] %3329;
                                                                                                                                                                                 u[2][223] = in_3[223] + e1[2][223] %3329;
                                                                                                                                                                                 u[2][224] = in_3[224] + e1[2][224] %3329;
                                                                                                                                                                                 u[2][225] = in_3[225] + e1[2][225] %3329;
                                                                                                                                                                                 u[2][226] = in_3[226] + e1[2][226] %3329;
                                                                                                                                                                                 u[2][227] = in_3[227] + e1[2][227] %3329;
                                                                                                                                                                                 u[2][228] = in_3[228] + e1[2][228] %3329;
                                                                                                                                                                                 u[2][229] = in_3[229] + e1[2][229] %3329;
                                                                                                                                                                                 u[2][230] = in_3[230] + e1[2][230] %3329;
                                                                                                                                                                                 u[2][231] = in_3[231] + e1[2][231] %3329;
                                                                                                                                                                                 u[2][232] = in_3[232] + e1[2][232] %3329;
                                                                                                                                                                                 u[2][233] = in_3[233] + e1[2][233] %3329;
                                                                                                                                                                                 u[2][234] = in_3[234] + e1[2][234] %3329;
                                                                                                                                                                                 u[2][235] = in_3[235] + e1[2][235] %3329;
                                                                                                                                                                                 u[2][236] = in_3[236] + e1[2][236] %3329;
                                                                                                                                                                                 u[2][237] = in_3[237] + e1[2][237] %3329;
                                                                                                                                                                                 u[2][238] = in_3[238] + e1[2][238] %3329;
                                                                                                                                                                                 u[2][239] = in_3[239] + e1[2][239] %3329;
                                                                                                                                                                                 u[2][240] = in_3[240] + e1[2][240] %3329;
                                                                                                                                                                                 u[2][241] = in_3[241] + e1[2][241] %3329;
                                                                                                                                                                                 u[2][242] = in_3[242] + e1[2][242] %3329;
                                                                                                                                                                                 u[2][243] = in_3[243] + e1[2][243] %3329;
                                                                                                                                                                                 u[2][244] = in_3[244] + e1[2][244] %3329;
                                                                                                                                                                                 u[2][245] = in_3[245] + e1[2][245] %3329;
                                                                                                                                                                                 u[2][246] = in_3[246] + e1[2][246] %3329;
                                                                                                                                                                                 u[2][247] = in_3[247] + e1[2][247] %3329;
                                                                                                                                                                                 u[2][248] = in_3[248] + e1[2][248] %3329;
                                                                                                                                                                                 u[2][249] = in_3[249] + e1[2][249] %3329;
                                                                                                                                                                                 u[2][250] = in_3[250] + e1[2][250] %3329;
                                                                                                                                                                                 u[2][251] = in_3[251] + e1[2][251] %3329;
                                                                                                                                                                                 u[2][252] = in_3[252] + e1[2][252] %3329;
                                                                                                                                                                                 u[2][253] = in_3[253] + e1[2][253] %3329;
                                                                                                                                                                                 u[2][254] = in_3[254] + e1[2][254] %3329;
                                                                                                                                                                                 u[2][255] = in_3[255] + e1[2][255] %3329;
                                                                                                                                                                                   v[0] = (in_4[0] + in_5[0] + in_6[0] + {16'b0, decom_out[0]} + {20'b0, e2[0]}) % 3329;
                                                                                                                                                                                     v[1] = (in_4[1] + in_5[1] + in_6[1] + {16'b0, decom_out[1]} + {20'b0, e2[1]}) % 3329;
                                                                                                                                                                                     v[2] = (in_4[2] + in_5[2] + in_6[2] + {16'b0, decom_out[2]} + {20'b0, e2[2]}) % 3329;
                                                                                                                                                                                     v[3] = (in_4[3] + in_5[3] + in_6[3] + {16'b0, decom_out[3]} + {20'b0, e2[3]}) % 3329;
                                                                                                                                                                                     v[4] = (in_4[4] + in_5[4] + in_6[4] + {16'b0, decom_out[4]} + {20'b0, e2[4]}) % 3329;
                                                                                                                                                                                     v[5] = (in_4[5] + in_5[5] + in_6[5] + {16'b0, decom_out[5]} + {20'b0, e2[5]}) % 3329;
                                                                                                                                                                                     v[6] = (in_4[6] + in_5[6] + in_6[6] + {16'b0, decom_out[6]} + {20'b0, e2[6]}) % 3329;
                                                                                                                                                                                     v[7] = (in_4[7] + in_5[7] + in_6[7] + {16'b0, decom_out[7]} + {20'b0, e2[7]}) % 3329;
                                                                                                                                                                                     v[8] = (in_4[8] + in_5[8] + in_6[8] + {16'b0, decom_out[8]} + {20'b0, e2[8]}) % 3329;
                                                                                                                                                                                     v[9] = (in_4[9] + in_5[9] + in_6[9] + {16'b0, decom_out[9]} + {20'b0, e2[9]}) % 3329;
                                                                                                                                                                                     v[10] = (in_4[10] + in_5[10] + in_6[10] + {16'b0, decom_out[10]} + {20'b0, e2[10]}) % 3329;
                                                                                                                                                                                     v[11] = (in_4[11] + in_5[11] + in_6[11] + {16'b0, decom_out[11]} + {20'b0, e2[11]}) % 3329;
                                                                                                                                                                                     v[12] = (in_4[12] + in_5[12] + in_6[12] + {16'b0, decom_out[12]} + {20'b0, e2[12]}) % 3329;
                                                                                                                                                                                     v[13] = (in_4[13] + in_5[13] + in_6[13] + {16'b0, decom_out[13]} + {20'b0, e2[13]}) % 3329;
                                                                                                                                                                                     v[14] = (in_4[14] + in_5[14] + in_6[14] + {16'b0, decom_out[14]} + {20'b0, e2[14]}) % 3329;
                                                                                                                                                                                     v[15] = (in_4[15] + in_5[15] + in_6[15] + {16'b0, decom_out[15]} + {20'b0, e2[15]}) % 3329;
                                                                                                                                                                                     v[16] = (in_4[16] + in_5[16] + in_6[16] + {16'b0, decom_out[16]} + {20'b0, e2[16]}) % 3329;
                                                                                                                                                                                     v[17] = (in_4[17] + in_5[17] + in_6[17] + {16'b0, decom_out[17]} + {20'b0, e2[17]}) % 3329;
                                                                                                                                                                                     v[18] = (in_4[18] + in_5[18] + in_6[18] + {16'b0, decom_out[18]} + {20'b0, e2[18]}) % 3329;
                                                                                                                                                                                     v[19] = (in_4[19] + in_5[19] + in_6[19] + {16'b0, decom_out[19]} + {20'b0, e2[19]}) % 3329;
                                                                                                                                                                                     v[20] = (in_4[20] + in_5[20] + in_6[20] + {16'b0, decom_out[20]} + {20'b0, e2[20]}) % 3329;
                                                                                                                                                                                     v[21] = (in_4[21] + in_5[21] + in_6[21] + {16'b0, decom_out[21]} + {20'b0, e2[21]}) % 3329;
                                                                                                                                                                                     v[22] = (in_4[22] + in_5[22] + in_6[22] + {16'b0, decom_out[22]} + {20'b0, e2[22]}) % 3329;
                                                                                                                                                                                     v[23] = (in_4[23] + in_5[23] + in_6[23] + {16'b0, decom_out[23]} + {20'b0, e2[23]}) % 3329;
                                                                                                                                                                                     v[24] = (in_4[24] + in_5[24] + in_6[24] + {16'b0, decom_out[24]} + {20'b0, e2[24]}) % 3329;
                                                                                                                                                                                     v[25] = (in_4[25] + in_5[25] + in_6[25] + {16'b0, decom_out[25]} + {20'b0, e2[25]}) % 3329;
                                                                                                                                                                                     v[26] = (in_4[26] + in_5[26] + in_6[26] + {16'b0, decom_out[26]} + {20'b0, e2[26]}) % 3329;
                                                                                                                                                                                     v[27] = (in_4[27] + in_5[27] + in_6[27] + {16'b0, decom_out[27]} + {20'b0, e2[27]}) % 3329;
                                                                                                                                                                                     v[28] = (in_4[28] + in_5[28] + in_6[28] + {16'b0, decom_out[28]} + {20'b0, e2[28]}) % 3329;
                                                                                                                                                                                     v[29] = (in_4[29] + in_5[29] + in_6[29] + {16'b0, decom_out[29]} + {20'b0, e2[29]}) % 3329;
                                                                                                                                                                                     v[30] = (in_4[30] + in_5[30] + in_6[30] + {16'b0, decom_out[30]} + {20'b0, e2[30]}) % 3329;
                                                                                                                                                                                     v[31] = (in_4[31] + in_5[31] + in_6[31] + {16'b0, decom_out[31]} + {20'b0, e2[31]}) % 3329;
                                                                                                                                                                                     v[32] = (in_4[32] + in_5[32] + in_6[32] + {16'b0, decom_out[32]} + {20'b0, e2[32]}) % 3329;
                                                                                                                                                                                     v[33] = (in_4[33] + in_5[33] + in_6[33] + {16'b0, decom_out[33]} + {20'b0, e2[33]}) % 3329;
                                                                                                                                                                                     v[34] = (in_4[34] + in_5[34] + in_6[34] + {16'b0, decom_out[34]} + {20'b0, e2[34]}) % 3329;
                                                                                                                                                                                     v[35] = (in_4[35] + in_5[35] + in_6[35] + {16'b0, decom_out[35]} + {20'b0, e2[35]}) % 3329;
                                                                                                                                                                                     v[36] = (in_4[36] + in_5[36] + in_6[36] + {16'b0, decom_out[36]} + {20'b0, e2[36]}) % 3329;
                                                                                                                                                                                     v[37] = (in_4[37] + in_5[37] + in_6[37] + {16'b0, decom_out[37]} + {20'b0, e2[37]}) % 3329;
                                                                                                                                                                                     v[38] = (in_4[38] + in_5[38] + in_6[38] + {16'b0, decom_out[38]} + {20'b0, e2[38]}) % 3329;
                                                                                                                                                                                     v[39] = (in_4[39] + in_5[39] + in_6[39] + {16'b0, decom_out[39]} + {20'b0, e2[39]}) % 3329;
                                                                                                                                                                                     v[40] = (in_4[40] + in_5[40] + in_6[40] + {16'b0, decom_out[40]} + {20'b0, e2[40]}) % 3329;
                                                                                                                                                                                     v[41] = (in_4[41] + in_5[41] + in_6[41] + {16'b0, decom_out[41]} + {20'b0, e2[41]}) % 3329;
                                                                                                                                                                                     v[42] = (in_4[42] + in_5[42] + in_6[42] + {16'b0, decom_out[42]} + {20'b0, e2[42]}) % 3329;
                                                                                                                                                                                     v[43] = (in_4[43] + in_5[43] + in_6[43] + {16'b0, decom_out[43]} + {20'b0, e2[43]}) % 3329;
                                                                                                                                                                                     v[44] = (in_4[44] + in_5[44] + in_6[44] + {16'b0, decom_out[44]} + {20'b0, e2[44]}) % 3329;
                                                                                                                                                                                     v[45] = (in_4[45] + in_5[45] + in_6[45] + {16'b0, decom_out[45]} + {20'b0, e2[45]}) % 3329;
                                                                                                                                                                                     v[46] = (in_4[46] + in_5[46] + in_6[46] + {16'b0, decom_out[46]} + {20'b0, e2[46]}) % 3329;
                                                                                                                                                                                     v[47] = (in_4[47] + in_5[47] + in_6[47] + {16'b0, decom_out[47]} + {20'b0, e2[47]}) % 3329;
                                                                                                                                                                                     v[48] = (in_4[48] + in_5[48] + in_6[48] + {16'b0, decom_out[48]} + {20'b0, e2[48]}) % 3329;
                                                                                                                                                                                     v[49] = (in_4[49] + in_5[49] + in_6[49] + {16'b0, decom_out[49]} + {20'b0, e2[49]}) % 3329;
                                                                                                                                                                                     v[50] = (in_4[50] + in_5[50] + in_6[50] + {16'b0, decom_out[50]} + {20'b0, e2[50]}) % 3329;
                                                                                                                                                                                     v[51] = (in_4[51] + in_5[51] + in_6[51] + {16'b0, decom_out[51]} + {20'b0, e2[51]}) % 3329;
                                                                                                                                                                                     v[52] = (in_4[52] + in_5[52] + in_6[52] + {16'b0, decom_out[52]} + {20'b0, e2[52]}) % 3329;
                                                                                                                                                                                     v[53] = (in_4[53] + in_5[53] + in_6[53] + {16'b0, decom_out[53]} + {20'b0, e2[53]}) % 3329;
                                                                                                                                                                                     v[54] = (in_4[54] + in_5[54] + in_6[54] + {16'b0, decom_out[54]} + {20'b0, e2[54]}) % 3329;
                                                                                                                                                                                     v[55] = (in_4[55] + in_5[55] + in_6[55] + {16'b0, decom_out[55]} + {20'b0, e2[55]}) % 3329;
                                                                                                                                                                                     v[56] = (in_4[56] + in_5[56] + in_6[56] + {16'b0, decom_out[56]} + {20'b0, e2[56]}) % 3329;
                                                                                                                                                                                     v[57] = (in_4[57] + in_5[57] + in_6[57] + {16'b0, decom_out[57]} + {20'b0, e2[57]}) % 3329;
                                                                                                                                                                                     v[58] = (in_4[58] + in_5[58] + in_6[58] + {16'b0, decom_out[58]} + {20'b0, e2[58]}) % 3329;
                                                                                                                                                                                     v[59] = (in_4[59] + in_5[59] + in_6[59] + {16'b0, decom_out[59]} + {20'b0, e2[59]}) % 3329;
                                                                                                                                                                                     v[60] = (in_4[60] + in_5[60] + in_6[60] + {16'b0, decom_out[60]} + {20'b0, e2[60]}) % 3329;
                                                                                                                                                                                     v[61] = (in_4[61] + in_5[61] + in_6[61] + {16'b0, decom_out[61]} + {20'b0, e2[61]}) % 3329;
                                                                                                                                                                                     v[62] = (in_4[62] + in_5[62] + in_6[62] + {16'b0, decom_out[62]} + {20'b0, e2[62]}) % 3329;
                                                                                                                                                                                     v[63] = (in_4[63] + in_5[63] + in_6[63] + {16'b0, decom_out[63]} + {20'b0, e2[63]}) % 3329;
                                                                                                                                                                                     v[64] = (in_4[64] + in_5[64] + in_6[64] + {16'b0, decom_out[64]} + {20'b0, e2[64]}) % 3329;
                                                                                                                                                                                     v[65] = (in_4[65] + in_5[65] + in_6[65] + {16'b0, decom_out[65]} + {20'b0, e2[65]}) % 3329;
                                                                                                                                                                                     v[66] = (in_4[66] + in_5[66] + in_6[66] + {16'b0, decom_out[66]} + {20'b0, e2[66]}) % 3329;
                                                                                                                                                                                     v[67] = (in_4[67] + in_5[67] + in_6[67] + {16'b0, decom_out[67]} + {20'b0, e2[67]}) % 3329;
                                                                                                                                                                                     v[68] = (in_4[68] + in_5[68] + in_6[68] + {16'b0, decom_out[68]} + {20'b0, e2[68]}) % 3329;
                                                                                                                                                                                     v[69] = (in_4[69] + in_5[69] + in_6[69] + {16'b0, decom_out[69]} + {20'b0, e2[69]}) % 3329;
                                                                                                                                                                                     v[70] = (in_4[70] + in_5[70] + in_6[70] + {16'b0, decom_out[70]} + {20'b0, e2[70]}) % 3329;
                                                                                                                                                                                     v[71] = (in_4[71] + in_5[71] + in_6[71] + {16'b0, decom_out[71]} + {20'b0, e2[71]}) % 3329;
                                                                                                                                                                                     v[72] = (in_4[72] + in_5[72] + in_6[72] + {16'b0, decom_out[72]} + {20'b0, e2[72]}) % 3329;
                                                                                                                                                                                     v[73] = (in_4[73] + in_5[73] + in_6[73] + {16'b0, decom_out[73]} + {20'b0, e2[73]}) % 3329;
                                                                                                                                                                                     v[74] = (in_4[74] + in_5[74] + in_6[74] + {16'b0, decom_out[74]} + {20'b0, e2[74]}) % 3329;
                                                                                                                                                                                     v[75] = (in_4[75] + in_5[75] + in_6[75] + {16'b0, decom_out[75]} + {20'b0, e2[75]}) % 3329;
                                                                                                                                                                                     v[76] = (in_4[76] + in_5[76] + in_6[76] + {16'b0, decom_out[76]} + {20'b0, e2[76]}) % 3329;
                                                                                                                                                                                     v[77] = (in_4[77] + in_5[77] + in_6[77] + {16'b0, decom_out[77]} + {20'b0, e2[77]}) % 3329;
                                                                                                                                                                                     v[78] = (in_4[78] + in_5[78] + in_6[78] + {16'b0, decom_out[78]} + {20'b0, e2[78]}) % 3329;
                                                                                                                                                                                     v[79] = (in_4[79] + in_5[79] + in_6[79] + {16'b0, decom_out[79]} + {20'b0, e2[79]}) % 3329;
                                                                                                                                                                                     v[80] = (in_4[80] + in_5[80] + in_6[80] + {16'b0, decom_out[80]} + {20'b0, e2[80]}) % 3329;
                                                                                                                                                                                     v[81] = (in_4[81] + in_5[81] + in_6[81] + {16'b0, decom_out[81]} + {20'b0, e2[81]}) % 3329;
                                                                                                                                                                                     v[82] = (in_4[82] + in_5[82] + in_6[82] + {16'b0, decom_out[82]} + {20'b0, e2[82]}) % 3329;
                                                                                                                                                                                     v[83] = (in_4[83] + in_5[83] + in_6[83] + {16'b0, decom_out[83]} + {20'b0, e2[83]}) % 3329;
                                                                                                                                                                                     v[84] = (in_4[84] + in_5[84] + in_6[84] + {16'b0, decom_out[84]} + {20'b0, e2[84]}) % 3329;
                                                                                                                                                                                     v[85] = (in_4[85] + in_5[85] + in_6[85] + {16'b0, decom_out[85]} + {20'b0, e2[85]}) % 3329;
                                                                                                                                                                                     v[86] = (in_4[86] + in_5[86] + in_6[86] + {16'b0, decom_out[86]} + {20'b0, e2[86]}) % 3329;
                                                                                                                                                                                     v[87] = (in_4[87] + in_5[87] + in_6[87] + {16'b0, decom_out[87]} + {20'b0, e2[87]}) % 3329;
                                                                                                                                                                                     v[88] = (in_4[88] + in_5[88] + in_6[88] + {16'b0, decom_out[88]} + {20'b0, e2[88]}) % 3329;
                                                                                                                                                                                     v[89] = (in_4[89] + in_5[89] + in_6[89] + {16'b0, decom_out[89]} + {20'b0, e2[89]}) % 3329;
                                                                                                                                                                                     v[90] = (in_4[90] + in_5[90] + in_6[90] + {16'b0, decom_out[90]} + {20'b0, e2[90]}) % 3329;
                                                                                                                                                                                     v[91] = (in_4[91] + in_5[91] + in_6[91] + {16'b0, decom_out[91]} + {20'b0, e2[91]}) % 3329;
                                                                                                                                                                                     v[92] = (in_4[92] + in_5[92] + in_6[92] + {16'b0, decom_out[92]} + {20'b0, e2[92]}) % 3329;
                                                                                                                                                                                     v[93] = (in_4[93] + in_5[93] + in_6[93] + {16'b0, decom_out[93]} + {20'b0, e2[93]}) % 3329;
                                                                                                                                                                                     v[94] = (in_4[94] + in_5[94] + in_6[94] + {16'b0, decom_out[94]} + {20'b0, e2[94]}) % 3329;
                                                                                                                                                                                     v[95] = (in_4[95] + in_5[95] + in_6[95] + {16'b0, decom_out[95]} + {20'b0, e2[95]}) % 3329;
                                                                                                                                                                                     v[96] = (in_4[96] + in_5[96] + in_6[96] + {16'b0, decom_out[96]} + {20'b0, e2[96]}) % 3329;
                                                                                                                                                                                     v[97] = (in_4[97] + in_5[97] + in_6[97] + {16'b0, decom_out[97]} + {20'b0, e2[97]}) % 3329;
                                                                                                                                                                                     v[98] = (in_4[98] + in_5[98] + in_6[98] + {16'b0, decom_out[98]} + {20'b0, e2[98]}) % 3329;
                                                                                                                                                                                     v[99] = (in_4[99] + in_5[99] + in_6[99] + {16'b0, decom_out[99]} + {20'b0, e2[99]}) % 3329;
                                                                                                                                                                                     v[100] = (in_4[100] + in_5[100] + in_6[100] + {16'b0, decom_out[100]} + {20'b0, e2[100]}) % 3329;
                                                                                                                                                                                     v[101] = (in_4[101] + in_5[101] + in_6[101] + {16'b0, decom_out[101]} + {20'b0, e2[101]}) % 3329;
                                                                                                                                                                                     v[102] = (in_4[102] + in_5[102] + in_6[102] + {16'b0, decom_out[102]} + {20'b0, e2[102]}) % 3329;
                                                                                                                                                                                     v[103] = (in_4[103] + in_5[103] + in_6[103] + {16'b0, decom_out[103]} + {20'b0, e2[103]}) % 3329;
                                                                                                                                                                                     v[104] = (in_4[104] + in_5[104] + in_6[104] + {16'b0, decom_out[104]} + {20'b0, e2[104]}) % 3329;
                                                                                                                                                                                     v[105] = (in_4[105] + in_5[105] + in_6[105] + {16'b0, decom_out[105]} + {20'b0, e2[105]}) % 3329;
                                                                                                                                                                                     v[106] = (in_4[106] + in_5[106] + in_6[106] + {16'b0, decom_out[106]} + {20'b0, e2[106]}) % 3329;
                                                                                                                                                                                     v[107] = (in_4[107] + in_5[107] + in_6[107] + {16'b0, decom_out[107]} + {20'b0, e2[107]}) % 3329;
                                                                                                                                                                                     v[108] = (in_4[108] + in_5[108] + in_6[108] + {16'b0, decom_out[108]} + {20'b0, e2[108]}) % 3329;
                                                                                                                                                                                     v[109] = (in_4[109] + in_5[109] + in_6[109] + {16'b0, decom_out[109]} + {20'b0, e2[109]}) % 3329;
                                                                                                                                                                                     v[110] = (in_4[110] + in_5[110] + in_6[110] + {16'b0, decom_out[110]} + {20'b0, e2[110]}) % 3329;
                                                                                                                                                                                     v[111] = (in_4[111] + in_5[111] + in_6[111] + {16'b0, decom_out[111]} + {20'b0, e2[111]}) % 3329;
                                                                                                                                                                                     v[112] = (in_4[112] + in_5[112] + in_6[112] + {16'b0, decom_out[112]} + {20'b0, e2[112]}) % 3329;
                                                                                                                                                                                     v[113] = (in_4[113] + in_5[113] + in_6[113] + {16'b0, decom_out[113]} + {20'b0, e2[113]}) % 3329;
                                                                                                                                                                                     v[114] = (in_4[114] + in_5[114] + in_6[114] + {16'b0, decom_out[114]} + {20'b0, e2[114]}) % 3329;
                                                                                                                                                                                     v[115] = (in_4[115] + in_5[115] + in_6[115] + {16'b0, decom_out[115]} + {20'b0, e2[115]}) % 3329;
                                                                                                                                                                                     v[116] = (in_4[116] + in_5[116] + in_6[116] + {16'b0, decom_out[116]} + {20'b0, e2[116]}) % 3329;
                                                                                                                                                                                     v[117] = (in_4[117] + in_5[117] + in_6[117] + {16'b0, decom_out[117]} + {20'b0, e2[117]}) % 3329;
                                                                                                                                                                                     v[118] = (in_4[118] + in_5[118] + in_6[118] + {16'b0, decom_out[118]} + {20'b0, e2[118]}) % 3329;
                                                                                                                                                                                     v[119] = (in_4[119] + in_5[119] + in_6[119] + {16'b0, decom_out[119]} + {20'b0, e2[119]}) % 3329;
                                                                                                                                                                                     v[120] = (in_4[120] + in_5[120] + in_6[120] + {16'b0, decom_out[120]} + {20'b0, e2[120]}) % 3329;
                                                                                                                                                                                     v[121] = (in_4[121] + in_5[121] + in_6[121] + {16'b0, decom_out[121]} + {20'b0, e2[121]}) % 3329;
                                                                                                                                                                                     v[122] = (in_4[122] + in_5[122] + in_6[122] + {16'b0, decom_out[122]} + {20'b0, e2[122]}) % 3329;
                                                                                                                                                                                     v[123] = (in_4[123] + in_5[123] + in_6[123] + {16'b0, decom_out[123]} + {20'b0, e2[123]}) % 3329;
                                                                                                                                                                                     v[124] = (in_4[124] + in_5[124] + in_6[124] + {16'b0, decom_out[124]} + {20'b0, e2[124]}) % 3329;
                                                                                                                                                                                     v[125] = (in_4[125] + in_5[125] + in_6[125] + {16'b0, decom_out[125]} + {20'b0, e2[125]}) % 3329;
                                                                                                                                                                                     v[126] = (in_4[126] + in_5[126] + in_6[126] + {16'b0, decom_out[126]} + {20'b0, e2[126]}) % 3329;
                                                                                                                                                                                     v[127] = (in_4[127] + in_5[127] + in_6[127] + {16'b0, decom_out[127]} + {20'b0, e2[127]}) % 3329;
                                                                                                                                                                                     v[128] = (in_4[128] + in_5[128] + in_6[128] + {16'b0, decom_out[128]} + {20'b0, e2[128]}) % 3329;
                                                                                                                                                                                     v[129] = (in_4[129] + in_5[129] + in_6[129] + {16'b0, decom_out[129]} + {20'b0, e2[129]}) % 3329;
                                                                                                                                                                                     v[130] = (in_4[130] + in_5[130] + in_6[130] + {16'b0, decom_out[130]} + {20'b0, e2[130]}) % 3329;
                                                                                                                                                                                     v[131] = (in_4[131] + in_5[131] + in_6[131] + {16'b0, decom_out[131]} + {20'b0, e2[131]}) % 3329;
                                                                                                                                                                                     v[132] = (in_4[132] + in_5[132] + in_6[132] + {16'b0, decom_out[132]} + {20'b0, e2[132]}) % 3329;
                                                                                                                                                                                     v[133] = (in_4[133] + in_5[133] + in_6[133] + {16'b0, decom_out[133]} + {20'b0, e2[133]}) % 3329;
                                                                                                                                                                                     v[134] = (in_4[134] + in_5[134] + in_6[134] + {16'b0, decom_out[134]} + {20'b0, e2[134]}) % 3329;
                                                                                                                                                                                     v[135] = (in_4[135] + in_5[135] + in_6[135] + {16'b0, decom_out[135]} + {20'b0, e2[135]}) % 3329;
                                                                                                                                                                                     v[136] = (in_4[136] + in_5[136] + in_6[136] + {16'b0, decom_out[136]} + {20'b0, e2[136]}) % 3329;
                                                                                                                                                                                     v[137] = (in_4[137] + in_5[137] + in_6[137] + {16'b0, decom_out[137]} + {20'b0, e2[137]}) % 3329;
                                                                                                                                                                                     v[138] = (in_4[138] + in_5[138] + in_6[138] + {16'b0, decom_out[138]} + {20'b0, e2[138]}) % 3329;
                                                                                                                                                                                     v[139] = (in_4[139] + in_5[139] + in_6[139] + {16'b0, decom_out[139]} + {20'b0, e2[139]}) % 3329;
                                                                                                                                                                                     v[140] = (in_4[140] + in_5[140] + in_6[140] + {16'b0, decom_out[140]} + {20'b0, e2[140]}) % 3329;
                                                                                                                                                                                     v[141] = (in_4[141] + in_5[141] + in_6[141] + {16'b0, decom_out[141]} + {20'b0, e2[141]}) % 3329;
                                                                                                                                                                                     v[142] = (in_4[142] + in_5[142] + in_6[142] + {16'b0, decom_out[142]} + {20'b0, e2[142]}) % 3329;
                                                                                                                                                                                     v[143] = (in_4[143] + in_5[143] + in_6[143] + {16'b0, decom_out[143]} + {20'b0, e2[143]}) % 3329;
                                                                                                                                                                                     v[144] = (in_4[144] + in_5[144] + in_6[144] + {16'b0, decom_out[144]} + {20'b0, e2[144]}) % 3329;
                                                                                                                                                                                     v[145] = (in_4[145] + in_5[145] + in_6[145] + {16'b0, decom_out[145]} + {20'b0, e2[145]}) % 3329;
                                                                                                                                                                                     v[146] = (in_4[146] + in_5[146] + in_6[146] + {16'b0, decom_out[146]} + {20'b0, e2[146]}) % 3329;
                                                                                                                                                                                     v[147] = (in_4[147] + in_5[147] + in_6[147] + {16'b0, decom_out[147]} + {20'b0, e2[147]}) % 3329;
                                                                                                                                                                                     v[148] = (in_4[148] + in_5[148] + in_6[148] + {16'b0, decom_out[148]} + {20'b0, e2[148]}) % 3329;
                                                                                                                                                                                     v[149] = (in_4[149] + in_5[149] + in_6[149] + {16'b0, decom_out[149]} + {20'b0, e2[149]}) % 3329;
                                                                                                                                                                                     v[150] = (in_4[150] + in_5[150] + in_6[150] + {16'b0, decom_out[150]} + {20'b0, e2[150]}) % 3329;
                                                                                                                                                                                     v[151] = (in_4[151] + in_5[151] + in_6[151] + {16'b0, decom_out[151]} + {20'b0, e2[151]}) % 3329;
                                                                                                                                                                                     v[152] = (in_4[152] + in_5[152] + in_6[152] + {16'b0, decom_out[152]} + {20'b0, e2[152]}) % 3329;
                                                                                                                                                                                     v[153] = (in_4[153] + in_5[153] + in_6[153] + {16'b0, decom_out[153]} + {20'b0, e2[153]}) % 3329;
                                                                                                                                                                                     v[154] = (in_4[154] + in_5[154] + in_6[154] + {16'b0, decom_out[154]} + {20'b0, e2[154]}) % 3329;
                                                                                                                                                                                     v[155] = (in_4[155] + in_5[155] + in_6[155] + {16'b0, decom_out[155]} + {20'b0, e2[155]}) % 3329;
                                                                                                                                                                                     v[156] = (in_4[156] + in_5[156] + in_6[156] + {16'b0, decom_out[156]} + {20'b0, e2[156]}) % 3329;
                                                                                                                                                                                     v[157] = (in_4[157] + in_5[157] + in_6[157] + {16'b0, decom_out[157]} + {20'b0, e2[157]}) % 3329;
                                                                                                                                                                                     v[158] = (in_4[158] + in_5[158] + in_6[158] + {16'b0, decom_out[158]} + {20'b0, e2[158]}) % 3329;
                                                                                                                                                                                     v[159] = (in_4[159] + in_5[159] + in_6[159] + {16'b0, decom_out[159]} + {20'b0, e2[159]}) % 3329;
                                                                                                                                                                                     v[160] = (in_4[160] + in_5[160] + in_6[160] + {16'b0, decom_out[160]} + {20'b0, e2[160]}) % 3329;
                                                                                                                                                                                     v[161] = (in_4[161] + in_5[161] + in_6[161] + {16'b0, decom_out[161]} + {20'b0, e2[161]}) % 3329;
                                                                                                                                                                                     v[162] = (in_4[162] + in_5[162] + in_6[162] + {16'b0, decom_out[162]} + {20'b0, e2[162]}) % 3329;
                                                                                                                                                                                     v[163] = (in_4[163] + in_5[163] + in_6[163] + {16'b0, decom_out[163]} + {20'b0, e2[163]}) % 3329;
                                                                                                                                                                                     v[164] = (in_4[164] + in_5[164] + in_6[164] + {16'b0, decom_out[164]} + {20'b0, e2[164]}) % 3329;
                                                                                                                                                                                     v[165] = (in_4[165] + in_5[165] + in_6[165] + {16'b0, decom_out[165]} + {20'b0, e2[165]}) % 3329;
                                                                                                                                                                                     v[166] = (in_4[166] + in_5[166] + in_6[166] + {16'b0, decom_out[166]} + {20'b0, e2[166]}) % 3329;
                                                                                                                                                                                     v[167] = (in_4[167] + in_5[167] + in_6[167] + {16'b0, decom_out[167]} + {20'b0, e2[167]}) % 3329;
                                                                                                                                                                                     v[168] = (in_4[168] + in_5[168] + in_6[168] + {16'b0, decom_out[168]} + {20'b0, e2[168]}) % 3329;
                                                                                                                                                                                     v[169] = (in_4[169] + in_5[169] + in_6[169] + {16'b0, decom_out[169]} + {20'b0, e2[169]}) % 3329;
                                                                                                                                                                                     v[170] = (in_4[170] + in_5[170] + in_6[170] + {16'b0, decom_out[170]} + {20'b0, e2[170]}) % 3329;
                                                                                                                                                                                     v[171] = (in_4[171] + in_5[171] + in_6[171] + {16'b0, decom_out[171]} + {20'b0, e2[171]}) % 3329;
                                                                                                                                                                                     v[172] = (in_4[172] + in_5[172] + in_6[172] + {16'b0, decom_out[172]} + {20'b0, e2[172]}) % 3329;
                                                                                                                                                                                     v[173] = (in_4[173] + in_5[173] + in_6[173] + {16'b0, decom_out[173]} + {20'b0, e2[173]}) % 3329;
                                                                                                                                                                                     v[174] = (in_4[174] + in_5[174] + in_6[174] + {16'b0, decom_out[174]} + {20'b0, e2[174]}) % 3329;
                                                                                                                                                                                     v[175] = (in_4[175] + in_5[175] + in_6[175] + {16'b0, decom_out[175]} + {20'b0, e2[175]}) % 3329;
                                                                                                                                                                                     v[176] = (in_4[176] + in_5[176] + in_6[176] + {16'b0, decom_out[176]} + {20'b0, e2[176]}) % 3329;
                                                                                                                                                                                     v[177] = (in_4[177] + in_5[177] + in_6[177] + {16'b0, decom_out[177]} + {20'b0, e2[177]}) % 3329;
                                                                                                                                                                                     v[178] = (in_4[178] + in_5[178] + in_6[178] + {16'b0, decom_out[178]} + {20'b0, e2[178]}) % 3329;
                                                                                                                                                                                     v[179] = (in_4[179] + in_5[179] + in_6[179] + {16'b0, decom_out[179]} + {20'b0, e2[179]}) % 3329;
                                                                                                                                                                                     v[180] = (in_4[180] + in_5[180] + in_6[180] + {16'b0, decom_out[180]} + {20'b0, e2[180]}) % 3329;
                                                                                                                                                                                     v[181] = (in_4[181] + in_5[181] + in_6[181] + {16'b0, decom_out[181]} + {20'b0, e2[181]}) % 3329;
                                                                                                                                                                                     v[182] = (in_4[182] + in_5[182] + in_6[182] + {16'b0, decom_out[182]} + {20'b0, e2[182]}) % 3329;
                                                                                                                                                                                     v[183] = (in_4[183] + in_5[183] + in_6[183] + {16'b0, decom_out[183]} + {20'b0, e2[183]}) % 3329;
                                                                                                                                                                                     v[184] = (in_4[184] + in_5[184] + in_6[184] + {16'b0, decom_out[184]} + {20'b0, e2[184]}) % 3329;
                                                                                                                                                                                     v[185] = (in_4[185] + in_5[185] + in_6[185] + {16'b0, decom_out[185]} + {20'b0, e2[185]}) % 3329;
                                                                                                                                                                                     v[186] = (in_4[186] + in_5[186] + in_6[186] + {16'b0, decom_out[186]} + {20'b0, e2[186]}) % 3329;
                                                                                                                                                                                     v[187] = (in_4[187] + in_5[187] + in_6[187] + {16'b0, decom_out[187]} + {20'b0, e2[187]}) % 3329;
                                                                                                                                                                                     v[188] = (in_4[188] + in_5[188] + in_6[188] + {16'b0, decom_out[188]} + {20'b0, e2[188]}) % 3329;
                                                                                                                                                                                     v[189] = (in_4[189] + in_5[189] + in_6[189] + {16'b0, decom_out[189]} + {20'b0, e2[189]}) % 3329;
                                                                                                                                                                                     v[190] = (in_4[190] + in_5[190] + in_6[190] + {16'b0, decom_out[190]} + {20'b0, e2[190]}) % 3329;
                                                                                                                                                                                     v[191] = (in_4[191] + in_5[191] + in_6[191] + {16'b0, decom_out[191]} + {20'b0, e2[191]}) % 3329;
                                                                                                                                                                                     v[192] = (in_4[192] + in_5[192] + in_6[192] + {16'b0, decom_out[192]} + {20'b0, e2[192]}) % 3329;
                                                                                                                                                                                     v[193] = (in_4[193] + in_5[193] + in_6[193] + {16'b0, decom_out[193]} + {20'b0, e2[193]}) % 3329;
                                                                                                                                                                                     v[194] = (in_4[194] + in_5[194] + in_6[194] + {16'b0, decom_out[194]} + {20'b0, e2[194]}) % 3329;
                                                                                                                                                                                     v[195] = (in_4[195] + in_5[195] + in_6[195] + {16'b0, decom_out[195]} + {20'b0, e2[195]}) % 3329;
                                                                                                                                                                                     v[196] = (in_4[196] + in_5[196] + in_6[196] + {16'b0, decom_out[196]} + {20'b0, e2[196]}) % 3329;
                                                                                                                                                                                     v[197] = (in_4[197] + in_5[197] + in_6[197] + {16'b0, decom_out[197]} + {20'b0, e2[197]}) % 3329;
                                                                                                                                                                                     v[198] = (in_4[198] + in_5[198] + in_6[198] + {16'b0, decom_out[198]} + {20'b0, e2[198]}) % 3329;
                                                                                                                                                                                     v[199] = (in_4[199] + in_5[199] + in_6[199] + {16'b0, decom_out[199]} + {20'b0, e2[199]}) % 3329;
                                                                                                                                                                                     v[200] = (in_4[200] + in_5[200] + in_6[200] + {16'b0, decom_out[200]} + {20'b0, e2[200]}) % 3329;
                                                                                                                                                                                     v[201] = (in_4[201] + in_5[201] + in_6[201] + {16'b0, decom_out[201]} + {20'b0, e2[201]}) % 3329;
                                                                                                                                                                                     v[202] = (in_4[202] + in_5[202] + in_6[202] + {16'b0, decom_out[202]} + {20'b0, e2[202]}) % 3329;
                                                                                                                                                                                     v[203] = (in_4[203] + in_5[203] + in_6[203] + {16'b0, decom_out[203]} + {20'b0, e2[203]}) % 3329;
                                                                                                                                                                                     v[204] = (in_4[204] + in_5[204] + in_6[204] + {16'b0, decom_out[204]} + {20'b0, e2[204]}) % 3329;
                                                                                                                                                                                     v[205] = (in_4[205] + in_5[205] + in_6[205] + {16'b0, decom_out[205]} + {20'b0, e2[205]}) % 3329;
                                                                                                                                                                                     v[206] = (in_4[206] + in_5[206] + in_6[206] + {16'b0, decom_out[206]} + {20'b0, e2[206]}) % 3329;
                                                                                                                                                                                     v[207] = (in_4[207] + in_5[207] + in_6[207] + {16'b0, decom_out[207]} + {20'b0, e2[207]}) % 3329;
                                                                                                                                                                                     v[208] = (in_4[208] + in_5[208] + in_6[208] + {16'b0, decom_out[208]} + {20'b0, e2[208]}) % 3329;
                                                                                                                                                                                     v[209] = (in_4[209] + in_5[209] + in_6[209] + {16'b0, decom_out[209]} + {20'b0, e2[209]}) % 3329;
                                                                                                                                                                                     v[210] = (in_4[210] + in_5[210] + in_6[210] + {16'b0, decom_out[210]} + {20'b0, e2[210]}) % 3329;
                                                                                                                                                                                     v[211] = (in_4[211] + in_5[211] + in_6[211] + {16'b0, decom_out[211]} + {20'b0, e2[211]}) % 3329;
                                                                                                                                                                                     v[212] = (in_4[212] + in_5[212] + in_6[212] + {16'b0, decom_out[212]} + {20'b0, e2[212]}) % 3329;
                                                                                                                                                                                     v[213] = (in_4[213] + in_5[213] + in_6[213] + {16'b0, decom_out[213]} + {20'b0, e2[213]}) % 3329;
                                                                                                                                                                                     v[214] = (in_4[214] + in_5[214] + in_6[214] + {16'b0, decom_out[214]} + {20'b0, e2[214]}) % 3329;
                                                                                                                                                                                     v[215] = (in_4[215] + in_5[215] + in_6[215] + {16'b0, decom_out[215]} + {20'b0, e2[215]}) % 3329;
                                                                                                                                                                                     v[216] = (in_4[216] + in_5[216] + in_6[216] + {16'b0, decom_out[216]} + {20'b0, e2[216]}) % 3329;
                                                                                                                                                                                     v[217] = (in_4[217] + in_5[217] + in_6[217] + {16'b0, decom_out[217]} + {20'b0, e2[217]}) % 3329;
                                                                                                                                                                                     v[218] = (in_4[218] + in_5[218] + in_6[218] + {16'b0, decom_out[218]} + {20'b0, e2[218]}) % 3329;
                                                                                                                                                                                     v[219] = (in_4[219] + in_5[219] + in_6[219] + {16'b0, decom_out[219]} + {20'b0, e2[219]}) % 3329;
                                                                                                                                                                                     v[220] = (in_4[220] + in_5[220] + in_6[220] + {16'b0, decom_out[220]} + {20'b0, e2[220]}) % 3329;
                                                                                                                                                                                     v[221] = (in_4[221] + in_5[221] + in_6[221] + {16'b0, decom_out[221]} + {20'b0, e2[221]}) % 3329;
                                                                                                                                                                                     v[222] = (in_4[222] + in_5[222] + in_6[222] + {16'b0, decom_out[222]} + {20'b0, e2[222]}) % 3329;
                                                                                                                                                                                     v[223] = (in_4[223] + in_5[223] + in_6[223] + {16'b0, decom_out[223]} + {20'b0, e2[223]}) % 3329;
                                                                                                                                                                                     v[224] = (in_4[224] + in_5[224] + in_6[224] + {16'b0, decom_out[224]} + {20'b0, e2[224]}) % 3329;
                                                                                                                                                                                     v[225] = (in_4[225] + in_5[225] + in_6[225] + {16'b0, decom_out[225]} + {20'b0, e2[225]}) % 3329;
                                                                                                                                                                                     v[226] = (in_4[226] + in_5[226] + in_6[226] + {16'b0, decom_out[226]} + {20'b0, e2[226]}) % 3329;
                                                                                                                                                                                     v[227] = (in_4[227] + in_5[227] + in_6[227] + {16'b0, decom_out[227]} + {20'b0, e2[227]}) % 3329;
                                                                                                                                                                                     v[228] = (in_4[228] + in_5[228] + in_6[228] + {16'b0, decom_out[228]} + {20'b0, e2[228]}) % 3329;
                                                                                                                                                                                     v[229] = (in_4[229] + in_5[229] + in_6[229] + {16'b0, decom_out[229]} + {20'b0, e2[229]}) % 3329;
                                                                                                                                                                                     v[230] = (in_4[230] + in_5[230] + in_6[230] + {16'b0, decom_out[230]} + {20'b0, e2[230]}) % 3329;
                                                                                                                                                                                     v[231] = (in_4[231] + in_5[231] + in_6[231] + {16'b0, decom_out[231]} + {20'b0, e2[231]}) % 3329;
                                                                                                                                                                                     v[232] = (in_4[232] + in_5[232] + in_6[232] + {16'b0, decom_out[232]} + {20'b0, e2[232]}) % 3329;
                                                                                                                                                                                     v[233] = (in_4[233] + in_5[233] + in_6[233] + {16'b0, decom_out[233]} + {20'b0, e2[233]}) % 3329;
                                                                                                                                                                                     v[234] = (in_4[234] + in_5[234] + in_6[234] + {16'b0, decom_out[234]} + {20'b0, e2[234]}) % 3329;
                                                                                                                                                                                     v[235] = (in_4[235] + in_5[235] + in_6[235] + {16'b0, decom_out[235]} + {20'b0, e2[235]}) % 3329;
                                                                                                                                                                                     v[236] = (in_4[236] + in_5[236] + in_6[236] + {16'b0, decom_out[236]} + {20'b0, e2[236]}) % 3329;
                                                                                                                                                                                     v[237] = (in_4[237] + in_5[237] + in_6[237] + {16'b0, decom_out[237]} + {20'b0, e2[237]}) % 3329;
                                                                                                                                                                                     v[238] = (in_4[238] + in_5[238] + in_6[238] + {16'b0, decom_out[238]} + {20'b0, e2[238]}) % 3329;
                                                                                                                                                                                     v[239] = (in_4[239] + in_5[239] + in_6[239] + {16'b0, decom_out[239]} + {20'b0, e2[239]}) % 3329;
                                                                                                                                                                                     v[240] = (in_4[240] + in_5[240] + in_6[240] + {16'b0, decom_out[240]} + {20'b0, e2[240]}) % 3329;
                                                                                                                                                                                     v[241] = (in_4[241] + in_5[241] + in_6[241] + {16'b0, decom_out[241]} + {20'b0, e2[241]}) % 3329;
                                                                                                                                                                                     v[242] = (in_4[242] + in_5[242] + in_6[242] + {16'b0, decom_out[242]} + {20'b0, e2[242]}) % 3329;
                                                                                                                                                                                     v[243] = (in_4[243] + in_5[243] + in_6[243] + {16'b0, decom_out[243]} + {20'b0, e2[243]}) % 3329;
                                                                                                                                                                                     v[244] = (in_4[244] + in_5[244] + in_6[244] + {16'b0, decom_out[244]} + {20'b0, e2[244]}) % 3329;
                                                                                                                                                                                     v[245] = (in_4[245] + in_5[245] + in_6[245] + {16'b0, decom_out[245]} + {20'b0, e2[245]}) % 3329;
                                                                                                                                                                                     v[246] = (in_4[246] + in_5[246] + in_6[246] + {16'b0, decom_out[246]} + {20'b0, e2[246]}) % 3329;
                                                                                                                                                                                     v[247] = (in_4[247] + in_5[247] + in_6[247] + {16'b0, decom_out[247]} + {20'b0, e2[247]}) % 3329;
                                                                                                                                                                                     v[248] = (in_4[248] + in_5[248] + in_6[248] + {16'b0, decom_out[248]} + {20'b0, e2[248]}) % 3329;
                                                                                                                                                                                     v[249] = (in_4[249] + in_5[249] + in_6[249] + {16'b0, decom_out[249]} + {20'b0, e2[249]}) % 3329;
                                                                                                                                                                                     v[250] = (in_4[250] + in_5[250] + in_6[250] + {16'b0, decom_out[250]} + {20'b0, e2[250]}) % 3329;
                                                                                                                                                                                     v[251] = (in_4[251] + in_5[251] + in_6[251] + {16'b0, decom_out[251]} + {20'b0, e2[251]}) % 3329;
                                                                                                                                                                                     v[252] = (in_4[252] + in_5[252] + in_6[252] + {16'b0, decom_out[252]} + {20'b0, e2[252]}) % 3329;
                                                                                                                                                                                     v[253] = (in_4[253] + in_5[253] + in_6[253] + {16'b0, decom_out[253]} + {20'b0, e2[253]}) % 3329;
                                                                                                                                                                                     v[254] = (in_4[254] + in_5[254] + in_6[254] + {16'b0, decom_out[254]} + {20'b0, e2[254]}) % 3329;
                                                                                                                                                                                     v[255] = (in_4[255] + in_5[255] + in_6[255] + {16'b0, decom_out[255]} + {20'b0, e2[255]}) % 3329;


                                                                                                                                                                                    
                                           
                                                                                                                                                  end
                                                                                                                                                  end
                                                                                                                                              
                                                                                                                                              
                                           
                                                                    
                                                      end
                                                      end       
                                       
                                    
                                   
                          endmodule